module demux_1x16(
    input a,
    input [3:0] sel,
    output reg [15:0] b
    );
    //reg [15:0] b;

    always @(*)
    begin
        case (sel)  //case statement with "sel"
            4'h0 : begin
                        b[0] = a;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h1 : begin
                        b[0] = 1'b0;
                        b[1] = a;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h2 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = a;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h3 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = a;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h4 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = a;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h5 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = a;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h6 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = a;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h7 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = a;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h8 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = a;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'h9 : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = a;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'ha : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = a;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'hb : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = a;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'hc : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = a;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'hd : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = a;
                        b[14] = 1'b0;
                        b[15] = 1'b0;
                   end
            4'he : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = a;
                        b[15] = 1'b0;
                   end
            4'hf : begin
                        b[0] = 1'b0;
                        b[1] = 1'b0;
                        b[2] = 1'b0;
                        b[3] = 1'b0;
                        b[4] = 1'b0;
                        b[5] = 1'b0;
                        b[6] = 1'b0;
                        b[7] = 1'b0;
                        b[8] = 1'b0;
                        b[9] = 1'b0;
                        b[10] = 1'b0;
                        b[11] = 1'b0;
                        b[12] = 1'b0;
                        b[13] = 1'b0;
                        b[14] = 1'b0;
                        b[15] = a;
                   end

        endcase
    end

endmodule
