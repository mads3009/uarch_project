module NOT (
   input a,
   output out
);

   nand2$ nand1 (out,a, a);
   
endmodule

