module ic_shifter_decode(clk,
                         rst_n,
                         w_fe_ld_buf,
                         w_icache_lower_data,
                         w_icache_upper_data,
                         r_icache_lower_data,
                         r_icache_upper_data,
                         w_EIP_to_use,
                         w_fe_ic_data_shifted,
                         w_pr_repne,
                         w_pr_cs_over,
                         w_pr_ss_over,
                         w_pr_ds_over,
                         w_pr_es_over,
                         w_pr_fs_over,
                         w_pr_gs_over,
                         w_pr_size_over,
                         w_pr_0f,
                         w_pr_pos,
                         w_mux_sel);



input  clk;
input  rst_n;
input  [1:0]  w_fe_ld_buf;
input  [127:0]w_icache_lower_data;
input  [127:0]w_icache_upper_data;
input  [127:0]r_icache_lower_data;
input  [127:0]r_icache_upper_data;
input  [31:0] w_EIP_to_use;
output [255:0]w_fe_ic_data_shifted;

output [3:0]  w_pr_repne;
output [3:0]  w_pr_cs_over;
output [3:0]  w_pr_ss_over;
output [3:0]  w_pr_ds_over;
output [3:0]  w_pr_es_over;
output [3:0]  w_pr_fs_over;
output [3:0]  w_pr_gs_over;
output [3:0]  w_pr_size_over;
output [3:0]  w_pr_0f;
output [3:0]  w_pr_pos;
output [2:0]  w_mux_sel;



register #128 u_icache_lower_data(.clk(clk), .rst_n(rst_n), .set_n(1'b1), .ld(w_fe_ld_buf[0]), .data_i(w_icache_lower_data), .data_o(r_icache_lower_data));
register #128 u_icache_upper_data(.clk(clk), .rst_n(rst_n), .set_n(1'b1), .ld(w_fe_ld_buf[1]), .data_i(w_icache_upper_data), .data_o(r_icache_upper_data));

wire [255:0]  w_ic_data_shifted_00;
wire [255:0]  w_ic_data_shifted_01;
wire [255:0]  w_ic_data_shifted_10;
wire [255:0]  w_ic_data_shifted_11;

//4 shifters
byte_rotate_right #32 u_ic_data_shifter_00(
  .amt(w_EIP_to_use[4:0]),
  .in({r_icache_upper_data, r_icache_lower_data}),
  .out(w_ic_data_shifted_00)
  );
byte_rotate_right #32 u_ic_data_shifter_01(
  .amt(w_EIP_to_use[4:0]),
  .in({r_icache_upper_data, w_icache_lower_data}),
  .out(w_ic_data_shifted_01)
  );
byte_rotate_right #32 u_ic_data_shifter_10(
  .amt(w_EIP_to_use[4:0]),
  .in({w_icache_upper_data, r_icache_lower_data}),
  .out(w_ic_data_shifted_10)
  );
byte_rotate_right #32 u_ic_data_shifter_11(
  .amt(w_EIP_to_use[4:0]),
  .in({w_icache_upper_data, w_icache_lower_data}),
  .out(w_ic_data_shifted_11)
  );

//Muxing between the shifters
mux_nbit_4x1 #256 u_w_fe_ic_data_shifted(.a0(w_ic_data_shifted_00), .a1(w_ic_data_shifted_01), .a2(w_ic_data_shifted_10), .a3(w_ic_data_shifted_11), .sel(w_fe_ld_buf), .out(w_fe_ic_data_shifted));

wire [511:0] c1c0;
wire [511:0] c1b0;
wire [511:0] b1c0;
wire [511:0] b1b0;


assign c1c0 = {w_icache_upper_data, w_icache_lower_data,w_icache_upper_data, w_icache_lower_data};
assign c1b0 = {w_icache_upper_data, r_icache_lower_data,w_icache_upper_data, r_icache_lower_data};
assign b1c0 = {r_icache_upper_data, w_icache_lower_data,r_icache_upper_data, w_icache_lower_data};
assign b1b0 = {r_icache_upper_data, r_icache_lower_data,r_icache_upper_data, r_icache_lower_data};


wire [2:0] w_mux_sel_c1c0_gen[31:0];
wire [2:0] w_mux_sel_c1b0_gen[31:0];
wire [2:0] w_mux_sel_b1c0_gen[31:0];
wire [2:0] w_mux_sel_b1b0_gen[31:0];

wire [2:0]w_mux_sel_c1c0;
wire [2:0]w_mux_sel_c1b0;
wire [2:0]w_mux_sel_b1c0;
wire [2:0]w_mux_sel_b1b0;

wire [3:0] w_pr_repne_c1c0_gen[31:0];
wire [3:0] w_pr_repne_c1b0_gen[31:0];
wire [3:0] w_pr_repne_b1c0_gen[31:0];
wire [3:0] w_pr_repne_b1b0_gen[31:0];

wire [3:0]w_pr_repne_c1c0;
wire [3:0]w_pr_repne_c1b0;
wire [3:0]w_pr_repne_b1c0;
wire [3:0]w_pr_repne_b1b0;


wire [3:0] w_pr_cs_over_c1c0_gen[31:0];
wire [3:0] w_pr_cs_over_c1b0_gen[31:0];
wire [3:0] w_pr_cs_over_b1c0_gen[31:0];
wire [3:0] w_pr_cs_over_b1b0_gen[31:0];

wire [3:0]w_pr_cs_over_c1c0;
wire [3:0]w_pr_cs_over_c1b0;
wire [3:0]w_pr_cs_over_b1c0;
wire [3:0]w_pr_cs_over_b1b0;

wire [3:0] w_pr_ss_over_c1c0_gen[31:0];
wire [3:0] w_pr_ss_over_c1b0_gen[31:0];
wire [3:0] w_pr_ss_over_b1c0_gen[31:0];
wire [3:0] w_pr_ss_over_b1b0_gen[31:0];

wire [3:0]w_pr_ss_over_c1c0;
wire [3:0]w_pr_ss_over_c1b0;
wire [3:0]w_pr_ss_over_b1c0;
wire [3:0]w_pr_ss_over_b1b0;

wire [3:0] w_pr_ds_over_c1c0_gen[31:0];
wire [3:0] w_pr_ds_over_c1b0_gen[31:0];
wire [3:0] w_pr_ds_over_b1c0_gen[31:0];
wire [3:0] w_pr_ds_over_b1b0_gen[31:0];

wire [3:0]w_pr_ds_over_c1c0;
wire [3:0]w_pr_ds_over_c1b0;
wire [3:0]w_pr_ds_over_b1c0;
wire [3:0]w_pr_ds_over_b1b0;

wire [3:0] w_pr_es_over_c1c0_gen[31:0];
wire [3:0] w_pr_es_over_c1b0_gen[31:0];
wire [3:0] w_pr_es_over_b1c0_gen[31:0];
wire [3:0] w_pr_es_over_b1b0_gen[31:0];

wire [3:0]w_pr_es_over_c1c0;
wire [3:0]w_pr_es_over_c1b0;
wire [3:0]w_pr_es_over_b1c0;
wire [3:0]w_pr_es_over_b1b0;

wire [3:0] w_pr_fs_over_c1c0_gen[31:0];
wire [3:0] w_pr_fs_over_c1b0_gen[31:0];
wire [3:0] w_pr_fs_over_b1c0_gen[31:0];
wire [3:0] w_pr_fs_over_b1b0_gen[31:0];

wire [3:0]w_pr_fs_over_c1c0;
wire [3:0]w_pr_fs_over_c1b0;
wire [3:0]w_pr_fs_over_b1c0;
wire [3:0]w_pr_fs_over_b1b0;

wire [3:0] w_pr_gs_over_c1c0_gen[31:0];
wire [3:0] w_pr_gs_over_c1b0_gen[31:0];
wire [3:0] w_pr_gs_over_b1c0_gen[31:0];
wire [3:0] w_pr_gs_over_b1b0_gen[31:0];

wire [3:0]w_pr_gs_over_c1c0;
wire [3:0]w_pr_gs_over_c1b0;
wire [3:0]w_pr_gs_over_b1c0;
wire [3:0]w_pr_gs_over_b1b0;

wire [3:0] w_pr_size_over_c1c0_gen[31:0];
wire [3:0] w_pr_size_over_c1b0_gen[31:0];
wire [3:0] w_pr_size_over_b1c0_gen[31:0];
wire [3:0] w_pr_size_over_b1b0_gen[31:0];

wire [3:0]w_pr_size_over_c1c0;
wire [3:0]w_pr_size_over_c1b0;
wire [3:0]w_pr_size_over_b1c0;
wire [3:0]w_pr_size_over_b1b0;

wire [3:0] w_pr_0f_c1c0_gen[31:0];
wire [3:0] w_pr_0f_c1b0_gen[31:0];
wire [3:0] w_pr_0f_b1c0_gen[31:0];
wire [3:0] w_pr_0f_b1b0_gen[31:0];

wire [3:0]w_pr_0f_c1c0;
wire [3:0]w_pr_0f_c1b0;
wire [3:0]w_pr_0f_b1c0;
wire [3:0]w_pr_0f_b1b0;

wire [3:0] w_pr_pos_c1c0_gen[31:0];
wire [3:0] w_pr_pos_c1b0_gen[31:0];
wire [3:0] w_pr_pos_b1c0_gen[31:0];
wire [3:0] w_pr_pos_b1b0_gen[31:0];

wire [3:0]w_pr_pos_c1c0;
wire [3:0]w_pr_pos_c1b0;
wire [3:0]w_pr_pos_b1c0;
wire [3:0]w_pr_pos_b1b0;

genvar i;
generate
  for (i=0; i<32; i=i+1) begin : fetch_dec1
fetch_to_decode u_fetch_decode1 (.de_lower_16bytes (        c1c0[((i*8)+31):i*8]), 
                                .w_pr_repne        (        w_pr_repne_c1c0_gen[i]),
                                .w_pr_cs_over      (      w_pr_cs_over_c1c0_gen[i]),
                                .w_pr_ss_over      (      w_pr_ss_over_c1c0_gen[i]),
                                .w_pr_ds_over      (      w_pr_ds_over_c1c0_gen[i]),
                                .w_pr_es_over      (      w_pr_es_over_c1c0_gen[i]),
                                .w_pr_fs_over      (      w_pr_fs_over_c1c0_gen[i]),
                                .w_pr_gs_over      (      w_pr_gs_over_c1c0_gen[i]),
                                .w_pr_size_over    (    w_pr_size_over_c1c0_gen[i]),
                                .w_pr_0f           (           w_pr_0f_c1c0_gen[i]),
                                .w_pr_pos          (          w_pr_pos_c1c0_gen[i]),
                                .w_mux_sel         (         w_mux_sel_c1c0_gen[i]));
  end
endgenerate

mux_nbit_32x1 #3 u_mux_sel1(.a0  (w_mux_sel_c1c0_gen[0 ]),  
                           .a1  (w_mux_sel_c1c0_gen[1 ]),
                           .a2  (w_mux_sel_c1c0_gen[2 ]),
                           .a3  (w_mux_sel_c1c0_gen[3 ]),
                           .a4  (w_mux_sel_c1c0_gen[4 ]),
                           .a5  (w_mux_sel_c1c0_gen[5 ]),
                           .a6  (w_mux_sel_c1c0_gen[6 ]),
                           .a7  (w_mux_sel_c1c0_gen[7 ]),
                           .a8  (w_mux_sel_c1c0_gen[8 ]),
                           .a9  (w_mux_sel_c1c0_gen[9 ]),
                           .a10 (w_mux_sel_c1c0_gen[10]),
                           .a11 (w_mux_sel_c1c0_gen[11]),
                           .a12 (w_mux_sel_c1c0_gen[12]),
                           .a13 (w_mux_sel_c1c0_gen[13]),
                           .a14 (w_mux_sel_c1c0_gen[14]),
                           .a15 (w_mux_sel_c1c0_gen[15]),
                           .a16 (w_mux_sel_c1c0_gen[16]),
                           .a17 (w_mux_sel_c1c0_gen[17]),
                           .a18 (w_mux_sel_c1c0_gen[18]),
                           .a19 (w_mux_sel_c1c0_gen[19]),
                           .a20 (w_mux_sel_c1c0_gen[20]),
                           .a21 (w_mux_sel_c1c0_gen[21]),
                           .a22 (w_mux_sel_c1c0_gen[22]),
                           .a23 (w_mux_sel_c1c0_gen[23]),
                           .a24 (w_mux_sel_c1c0_gen[24]),
                           .a25 (w_mux_sel_c1c0_gen[25]),
                           .a26 (w_mux_sel_c1c0_gen[26]),
                           .a27 (w_mux_sel_c1c0_gen[27]),
                           .a28 (w_mux_sel_c1c0_gen[28]),
                           .a29 (w_mux_sel_c1c0_gen[29]),
                           .a30 (w_mux_sel_c1c0_gen[30]),
                           .a31 (w_mux_sel_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_mux_sel_c1c0));


mux_nbit_32x1 #4 u_pr_repn1(.a0  (w_pr_repne_c1c0_gen[0 ]),  
                           .a1  (w_pr_repne_c1c0_gen[1 ]),
                           .a2  (w_pr_repne_c1c0_gen[2 ]),
                           .a3  (w_pr_repne_c1c0_gen[3 ]),
                           .a4  (w_pr_repne_c1c0_gen[4 ]),
                           .a5  (w_pr_repne_c1c0_gen[5 ]),
                           .a6  (w_pr_repne_c1c0_gen[6 ]),
                           .a7  (w_pr_repne_c1c0_gen[7 ]),
                           .a8  (w_pr_repne_c1c0_gen[8 ]),
                           .a9  (w_pr_repne_c1c0_gen[9 ]),
                           .a10 (w_pr_repne_c1c0_gen[10]),
                           .a11 (w_pr_repne_c1c0_gen[11]),
                           .a12 (w_pr_repne_c1c0_gen[12]),
                           .a13 (w_pr_repne_c1c0_gen[13]),
                           .a14 (w_pr_repne_c1c0_gen[14]),
                           .a15 (w_pr_repne_c1c0_gen[15]),
                           .a16 (w_pr_repne_c1c0_gen[16]),
                           .a17 (w_pr_repne_c1c0_gen[17]),
                           .a18 (w_pr_repne_c1c0_gen[18]),
                           .a19 (w_pr_repne_c1c0_gen[19]),
                           .a20 (w_pr_repne_c1c0_gen[20]),
                           .a21 (w_pr_repne_c1c0_gen[21]),
                           .a22 (w_pr_repne_c1c0_gen[22]),
                           .a23 (w_pr_repne_c1c0_gen[23]),
                           .a24 (w_pr_repne_c1c0_gen[24]),
                           .a25 (w_pr_repne_c1c0_gen[25]),
                           .a26 (w_pr_repne_c1c0_gen[26]),
                           .a27 (w_pr_repne_c1c0_gen[27]),
                           .a28 (w_pr_repne_c1c0_gen[28]),
                           .a29 (w_pr_repne_c1c0_gen[29]),
                           .a30 (w_pr_repne_c1c0_gen[30]),
                           .a31 (w_pr_repne_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_repne_c1c0));


mux_nbit_32x1 #4 u_pr_cs1  (.a0  (w_pr_cs_over_c1c0_gen[0 ]),  
                           .a1  (w_pr_cs_over_c1c0_gen[1 ]),
                           .a2  (w_pr_cs_over_c1c0_gen[2 ]),
                           .a3  (w_pr_cs_over_c1c0_gen[3 ]),
                           .a4  (w_pr_cs_over_c1c0_gen[4 ]),
                           .a5  (w_pr_cs_over_c1c0_gen[5 ]),
                           .a6  (w_pr_cs_over_c1c0_gen[6 ]),
                           .a7  (w_pr_cs_over_c1c0_gen[7 ]),
                           .a8  (w_pr_cs_over_c1c0_gen[8 ]),
                           .a9  (w_pr_cs_over_c1c0_gen[9 ]),
                           .a10 (w_pr_cs_over_c1c0_gen[10]),
                           .a11 (w_pr_cs_over_c1c0_gen[11]),
                           .a12 (w_pr_cs_over_c1c0_gen[12]),
                           .a13 (w_pr_cs_over_c1c0_gen[13]),
                           .a14 (w_pr_cs_over_c1c0_gen[14]),
                           .a15 (w_pr_cs_over_c1c0_gen[15]),
                           .a16 (w_pr_cs_over_c1c0_gen[16]),
                           .a17 (w_pr_cs_over_c1c0_gen[17]),
                           .a18 (w_pr_cs_over_c1c0_gen[18]),
                           .a19 (w_pr_cs_over_c1c0_gen[19]),
                           .a20 (w_pr_cs_over_c1c0_gen[20]),
                           .a21 (w_pr_cs_over_c1c0_gen[21]),
                           .a22 (w_pr_cs_over_c1c0_gen[22]),
                           .a23 (w_pr_cs_over_c1c0_gen[23]),
                           .a24 (w_pr_cs_over_c1c0_gen[24]),
                           .a25 (w_pr_cs_over_c1c0_gen[25]),
                           .a26 (w_pr_cs_over_c1c0_gen[26]),
                           .a27 (w_pr_cs_over_c1c0_gen[27]),
                           .a28 (w_pr_cs_over_c1c0_gen[28]),
                           .a29 (w_pr_cs_over_c1c0_gen[29]),
                           .a30 (w_pr_cs_over_c1c0_gen[30]),
                           .a31 (w_pr_cs_over_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_cs_over_c1c0));

mux_nbit_32x1 #4 u_pr_ss1  (.a0  (w_pr_ss_over_c1c0_gen[0 ]),  
                           .a1  (w_pr_ss_over_c1c0_gen[1 ]),
                           .a2  (w_pr_ss_over_c1c0_gen[2 ]),
                           .a3  (w_pr_ss_over_c1c0_gen[3 ]),
                           .a4  (w_pr_ss_over_c1c0_gen[4 ]),
                           .a5  (w_pr_ss_over_c1c0_gen[5 ]),
                           .a6  (w_pr_ss_over_c1c0_gen[6 ]),
                           .a7  (w_pr_ss_over_c1c0_gen[7 ]),
                           .a8  (w_pr_ss_over_c1c0_gen[8 ]),
                           .a9  (w_pr_ss_over_c1c0_gen[9 ]),
                           .a10 (w_pr_ss_over_c1c0_gen[10]),
                           .a11 (w_pr_ss_over_c1c0_gen[11]),
                           .a12 (w_pr_ss_over_c1c0_gen[12]),
                           .a13 (w_pr_ss_over_c1c0_gen[13]),
                           .a14 (w_pr_ss_over_c1c0_gen[14]),
                           .a15 (w_pr_ss_over_c1c0_gen[15]),
                           .a16 (w_pr_ss_over_c1c0_gen[16]),
                           .a17 (w_pr_ss_over_c1c0_gen[17]),
                           .a18 (w_pr_ss_over_c1c0_gen[18]),
                           .a19 (w_pr_ss_over_c1c0_gen[19]),
                           .a20 (w_pr_ss_over_c1c0_gen[20]),
                           .a21 (w_pr_ss_over_c1c0_gen[21]),
                           .a22 (w_pr_ss_over_c1c0_gen[22]),
                           .a23 (w_pr_ss_over_c1c0_gen[23]),
                           .a24 (w_pr_ss_over_c1c0_gen[24]),
                           .a25 (w_pr_ss_over_c1c0_gen[25]),
                           .a26 (w_pr_ss_over_c1c0_gen[26]),
                           .a27 (w_pr_ss_over_c1c0_gen[27]),
                           .a28 (w_pr_ss_over_c1c0_gen[28]),
                           .a29 (w_pr_ss_over_c1c0_gen[29]),
                           .a30 (w_pr_ss_over_c1c0_gen[30]),
                           .a31 (w_pr_ss_over_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ss_over_c1c0));

mux_nbit_32x1 #4 u_pr_ds1  (.a0  (w_pr_ds_over_c1c0_gen[0 ]),  
                           .a1  (w_pr_ds_over_c1c0_gen[1 ]),
                           .a2  (w_pr_ds_over_c1c0_gen[2 ]),
                           .a3  (w_pr_ds_over_c1c0_gen[3 ]),
                           .a4  (w_pr_ds_over_c1c0_gen[4 ]),
                           .a5  (w_pr_ds_over_c1c0_gen[5 ]),
                           .a6  (w_pr_ds_over_c1c0_gen[6 ]),
                           .a7  (w_pr_ds_over_c1c0_gen[7 ]),
                           .a8  (w_pr_ds_over_c1c0_gen[8 ]),
                           .a9  (w_pr_ds_over_c1c0_gen[9 ]),
                           .a10 (w_pr_ds_over_c1c0_gen[10]),
                           .a11 (w_pr_ds_over_c1c0_gen[11]),
                           .a12 (w_pr_ds_over_c1c0_gen[12]),
                           .a13 (w_pr_ds_over_c1c0_gen[13]),
                           .a14 (w_pr_ds_over_c1c0_gen[14]),
                           .a15 (w_pr_ds_over_c1c0_gen[15]),
                           .a16 (w_pr_ds_over_c1c0_gen[16]),
                           .a17 (w_pr_ds_over_c1c0_gen[17]),
                           .a18 (w_pr_ds_over_c1c0_gen[18]),
                           .a19 (w_pr_ds_over_c1c0_gen[19]),
                           .a20 (w_pr_ds_over_c1c0_gen[20]),
                           .a21 (w_pr_ds_over_c1c0_gen[21]),
                           .a22 (w_pr_ds_over_c1c0_gen[22]),
                           .a23 (w_pr_ds_over_c1c0_gen[23]),
                           .a24 (w_pr_ds_over_c1c0_gen[24]),
                           .a25 (w_pr_ds_over_c1c0_gen[25]),
                           .a26 (w_pr_ds_over_c1c0_gen[26]),
                           .a27 (w_pr_ds_over_c1c0_gen[27]),
                           .a28 (w_pr_ds_over_c1c0_gen[28]),
                           .a29 (w_pr_ds_over_c1c0_gen[29]),
                           .a30 (w_pr_ds_over_c1c0_gen[30]),
                           .a31 (w_pr_ds_over_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ds_over_c1c0));

mux_nbit_32x1 #4 u_pr_es1  (.a0  (w_pr_es_over_c1c0_gen[0 ]),  
                           .a1  (w_pr_es_over_c1c0_gen[1 ]),
                           .a2  (w_pr_es_over_c1c0_gen[2 ]),
                           .a3  (w_pr_es_over_c1c0_gen[3 ]),
                           .a4  (w_pr_es_over_c1c0_gen[4 ]),
                           .a5  (w_pr_es_over_c1c0_gen[5 ]),
                           .a6  (w_pr_es_over_c1c0_gen[6 ]),
                           .a7  (w_pr_es_over_c1c0_gen[7 ]),
                           .a8  (w_pr_es_over_c1c0_gen[8 ]),
                           .a9  (w_pr_es_over_c1c0_gen[9 ]),
                           .a10 (w_pr_es_over_c1c0_gen[10]),
                           .a11 (w_pr_es_over_c1c0_gen[11]),
                           .a12 (w_pr_es_over_c1c0_gen[12]),
                           .a13 (w_pr_es_over_c1c0_gen[13]),
                           .a14 (w_pr_es_over_c1c0_gen[14]),
                           .a15 (w_pr_es_over_c1c0_gen[15]),
                           .a16 (w_pr_es_over_c1c0_gen[16]),
                           .a17 (w_pr_es_over_c1c0_gen[17]),
                           .a18 (w_pr_es_over_c1c0_gen[18]),
                           .a19 (w_pr_es_over_c1c0_gen[19]),
                           .a20 (w_pr_es_over_c1c0_gen[20]),
                           .a21 (w_pr_es_over_c1c0_gen[21]),
                           .a22 (w_pr_es_over_c1c0_gen[22]),
                           .a23 (w_pr_es_over_c1c0_gen[23]),
                           .a24 (w_pr_es_over_c1c0_gen[24]),
                           .a25 (w_pr_es_over_c1c0_gen[25]),
                           .a26 (w_pr_es_over_c1c0_gen[26]),
                           .a27 (w_pr_es_over_c1c0_gen[27]),
                           .a28 (w_pr_es_over_c1c0_gen[28]),
                           .a29 (w_pr_es_over_c1c0_gen[29]),
                           .a30 (w_pr_es_over_c1c0_gen[30]),
                           .a31 (w_pr_es_over_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_es_over_c1c0));

mux_nbit_32x1 #4 u_pr_fs1  (.a0  (w_pr_fs_over_c1c0_gen[0 ]),  
                           .a1  (w_pr_fs_over_c1c0_gen[1 ]),
                           .a2  (w_pr_fs_over_c1c0_gen[2 ]),
                           .a3  (w_pr_fs_over_c1c0_gen[3 ]),
                           .a4  (w_pr_fs_over_c1c0_gen[4 ]),
                           .a5  (w_pr_fs_over_c1c0_gen[5 ]),
                           .a6  (w_pr_fs_over_c1c0_gen[6 ]),
                           .a7  (w_pr_fs_over_c1c0_gen[7 ]),
                           .a8  (w_pr_fs_over_c1c0_gen[8 ]),
                           .a9  (w_pr_fs_over_c1c0_gen[9 ]),
                           .a10 (w_pr_fs_over_c1c0_gen[10]),
                           .a11 (w_pr_fs_over_c1c0_gen[11]),
                           .a12 (w_pr_fs_over_c1c0_gen[12]),
                           .a13 (w_pr_fs_over_c1c0_gen[13]),
                           .a14 (w_pr_fs_over_c1c0_gen[14]),
                           .a15 (w_pr_fs_over_c1c0_gen[15]),
                           .a16 (w_pr_fs_over_c1c0_gen[16]),
                           .a17 (w_pr_fs_over_c1c0_gen[17]),
                           .a18 (w_pr_fs_over_c1c0_gen[18]),
                           .a19 (w_pr_fs_over_c1c0_gen[19]),
                           .a20 (w_pr_fs_over_c1c0_gen[20]),
                           .a21 (w_pr_fs_over_c1c0_gen[21]),
                           .a22 (w_pr_fs_over_c1c0_gen[22]),
                           .a23 (w_pr_fs_over_c1c0_gen[23]),
                           .a24 (w_pr_fs_over_c1c0_gen[24]),
                           .a25 (w_pr_fs_over_c1c0_gen[25]),
                           .a26 (w_pr_fs_over_c1c0_gen[26]),
                           .a27 (w_pr_fs_over_c1c0_gen[27]),
                           .a28 (w_pr_fs_over_c1c0_gen[28]),
                           .a29 (w_pr_fs_over_c1c0_gen[29]),
                           .a30 (w_pr_fs_over_c1c0_gen[30]),
                           .a31 (w_pr_fs_over_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_fs_over_c1c0));

mux_nbit_32x1 #4 u_pr_gs1  (.a0  (w_pr_gs_over_c1c0_gen[0 ]),  
                           .a1  (w_pr_gs_over_c1c0_gen[1 ]),
                           .a2  (w_pr_gs_over_c1c0_gen[2 ]),
                           .a3  (w_pr_gs_over_c1c0_gen[3 ]),
                           .a4  (w_pr_gs_over_c1c0_gen[4 ]),
                           .a5  (w_pr_gs_over_c1c0_gen[5 ]),
                           .a6  (w_pr_gs_over_c1c0_gen[6 ]),
                           .a7  (w_pr_gs_over_c1c0_gen[7 ]),
                           .a8  (w_pr_gs_over_c1c0_gen[8 ]),
                           .a9  (w_pr_gs_over_c1c0_gen[9 ]),
                           .a10 (w_pr_gs_over_c1c0_gen[10]),
                           .a11 (w_pr_gs_over_c1c0_gen[11]),
                           .a12 (w_pr_gs_over_c1c0_gen[12]),
                           .a13 (w_pr_gs_over_c1c0_gen[13]),
                           .a14 (w_pr_gs_over_c1c0_gen[14]),
                           .a15 (w_pr_gs_over_c1c0_gen[15]),
                           .a16 (w_pr_gs_over_c1c0_gen[16]),
                           .a17 (w_pr_gs_over_c1c0_gen[17]),
                           .a18 (w_pr_gs_over_c1c0_gen[18]),
                           .a19 (w_pr_gs_over_c1c0_gen[19]),
                           .a20 (w_pr_gs_over_c1c0_gen[20]),
                           .a21 (w_pr_gs_over_c1c0_gen[21]),
                           .a22 (w_pr_gs_over_c1c0_gen[22]),
                           .a23 (w_pr_gs_over_c1c0_gen[23]),
                           .a24 (w_pr_gs_over_c1c0_gen[24]),
                           .a25 (w_pr_gs_over_c1c0_gen[25]),
                           .a26 (w_pr_gs_over_c1c0_gen[26]),
                           .a27 (w_pr_gs_over_c1c0_gen[27]),
                           .a28 (w_pr_gs_over_c1c0_gen[28]),
                           .a29 (w_pr_gs_over_c1c0_gen[29]),
                           .a30 (w_pr_gs_over_c1c0_gen[30]),
                           .a31 (w_pr_gs_over_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_gs_over_c1c0));

mux_nbit_32x1 #4 u_pr_size1(.a0  (w_pr_size_over_c1c0_gen[0 ]),  
                           .a1  (w_pr_size_over_c1c0_gen[1 ]),
                           .a2  (w_pr_size_over_c1c0_gen[2 ]),
                           .a3  (w_pr_size_over_c1c0_gen[3 ]),
                           .a4  (w_pr_size_over_c1c0_gen[4 ]),
                           .a5  (w_pr_size_over_c1c0_gen[5 ]),
                           .a6  (w_pr_size_over_c1c0_gen[6 ]),
                           .a7  (w_pr_size_over_c1c0_gen[7 ]),
                           .a8  (w_pr_size_over_c1c0_gen[8 ]),
                           .a9  (w_pr_size_over_c1c0_gen[9 ]),
                           .a10 (w_pr_size_over_c1c0_gen[10]),
                           .a11 (w_pr_size_over_c1c0_gen[11]),
                           .a12 (w_pr_size_over_c1c0_gen[12]),
                           .a13 (w_pr_size_over_c1c0_gen[13]),
                           .a14 (w_pr_size_over_c1c0_gen[14]),
                           .a15 (w_pr_size_over_c1c0_gen[15]),
                           .a16 (w_pr_size_over_c1c0_gen[16]),
                           .a17 (w_pr_size_over_c1c0_gen[17]),
                           .a18 (w_pr_size_over_c1c0_gen[18]),
                           .a19 (w_pr_size_over_c1c0_gen[19]),
                           .a20 (w_pr_size_over_c1c0_gen[20]),
                           .a21 (w_pr_size_over_c1c0_gen[21]),
                           .a22 (w_pr_size_over_c1c0_gen[22]),
                           .a23 (w_pr_size_over_c1c0_gen[23]),
                           .a24 (w_pr_size_over_c1c0_gen[24]),
                           .a25 (w_pr_size_over_c1c0_gen[25]),
                           .a26 (w_pr_size_over_c1c0_gen[26]),
                           .a27 (w_pr_size_over_c1c0_gen[27]),
                           .a28 (w_pr_size_over_c1c0_gen[28]),
                           .a29 (w_pr_size_over_c1c0_gen[29]),
                           .a30 (w_pr_size_over_c1c0_gen[30]),
                           .a31 (w_pr_size_over_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_size_over_c1c0));

mux_nbit_32x1 #4 u_pr_0f1  (.a0  (w_pr_0f_c1c0_gen[0 ]),  
                           .a1  (w_pr_0f_c1c0_gen[1 ]),
                           .a2  (w_pr_0f_c1c0_gen[2 ]),
                           .a3  (w_pr_0f_c1c0_gen[3 ]),
                           .a4  (w_pr_0f_c1c0_gen[4 ]),
                           .a5  (w_pr_0f_c1c0_gen[5 ]),
                           .a6  (w_pr_0f_c1c0_gen[6 ]),
                           .a7  (w_pr_0f_c1c0_gen[7 ]),
                           .a8  (w_pr_0f_c1c0_gen[8 ]),
                           .a9  (w_pr_0f_c1c0_gen[9 ]),
                           .a10 (w_pr_0f_c1c0_gen[10]),
                           .a11 (w_pr_0f_c1c0_gen[11]),
                           .a12 (w_pr_0f_c1c0_gen[12]),
                           .a13 (w_pr_0f_c1c0_gen[13]),
                           .a14 (w_pr_0f_c1c0_gen[14]),
                           .a15 (w_pr_0f_c1c0_gen[15]),
                           .a16 (w_pr_0f_c1c0_gen[16]),
                           .a17 (w_pr_0f_c1c0_gen[17]),
                           .a18 (w_pr_0f_c1c0_gen[18]),
                           .a19 (w_pr_0f_c1c0_gen[19]),
                           .a20 (w_pr_0f_c1c0_gen[20]),
                           .a21 (w_pr_0f_c1c0_gen[21]),
                           .a22 (w_pr_0f_c1c0_gen[22]),
                           .a23 (w_pr_0f_c1c0_gen[23]),
                           .a24 (w_pr_0f_c1c0_gen[24]),
                           .a25 (w_pr_0f_c1c0_gen[25]),
                           .a26 (w_pr_0f_c1c0_gen[26]),
                           .a27 (w_pr_0f_c1c0_gen[27]),
                           .a28 (w_pr_0f_c1c0_gen[28]),
                           .a29 (w_pr_0f_c1c0_gen[29]),
                           .a30 (w_pr_0f_c1c0_gen[30]),
                           .a31 (w_pr_0f_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_0f_c1c0));

mux_nbit_32x1 #4 u_pr_pos1  (.a0  (w_pr_pos_c1c0_gen[0 ]),  
                           .a1  (w_pr_pos_c1c0_gen[1 ]),
                           .a2  (w_pr_pos_c1c0_gen[2 ]),
                           .a3  (w_pr_pos_c1c0_gen[3 ]),
                           .a4  (w_pr_pos_c1c0_gen[4 ]),
                           .a5  (w_pr_pos_c1c0_gen[5 ]),
                           .a6  (w_pr_pos_c1c0_gen[6 ]),
                           .a7  (w_pr_pos_c1c0_gen[7 ]),
                           .a8  (w_pr_pos_c1c0_gen[8 ]),
                           .a9  (w_pr_pos_c1c0_gen[9 ]),
                           .a10 (w_pr_pos_c1c0_gen[10]),
                           .a11 (w_pr_pos_c1c0_gen[11]),
                           .a12 (w_pr_pos_c1c0_gen[12]),
                           .a13 (w_pr_pos_c1c0_gen[13]),
                           .a14 (w_pr_pos_c1c0_gen[14]),
                           .a15 (w_pr_pos_c1c0_gen[15]),
                           .a16 (w_pr_pos_c1c0_gen[16]),
                           .a17 (w_pr_pos_c1c0_gen[17]),
                           .a18 (w_pr_pos_c1c0_gen[18]),
                           .a19 (w_pr_pos_c1c0_gen[19]),
                           .a20 (w_pr_pos_c1c0_gen[20]),
                           .a21 (w_pr_pos_c1c0_gen[21]),
                           .a22 (w_pr_pos_c1c0_gen[22]),
                           .a23 (w_pr_pos_c1c0_gen[23]),
                           .a24 (w_pr_pos_c1c0_gen[24]),
                           .a25 (w_pr_pos_c1c0_gen[25]),
                           .a26 (w_pr_pos_c1c0_gen[26]),
                           .a27 (w_pr_pos_c1c0_gen[27]),
                           .a28 (w_pr_pos_c1c0_gen[28]),
                           .a29 (w_pr_pos_c1c0_gen[29]),
                           .a30 (w_pr_pos_c1c0_gen[30]),
                           .a31 (w_pr_pos_c1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_pos_c1c0));


//c1b0

generate
  for (i=0; i<32; i=i+1) begin : fetch_dec2
fetch_to_decode u_fetch_decode2 (.de_lower_16bytes  (        c1b0[((i*8)+31):i*8]), 
                                .w_pr_repne        (        w_pr_repne_c1b0_gen[i]),
                                .w_pr_cs_over      (      w_pr_cs_over_c1b0_gen[i]),
                                .w_pr_ss_over      (      w_pr_ss_over_c1b0_gen[i]),
                                .w_pr_ds_over      (      w_pr_ds_over_c1b0_gen[i]),
                                .w_pr_es_over      (      w_pr_es_over_c1b0_gen[i]),
                                .w_pr_fs_over      (      w_pr_fs_over_c1b0_gen[i]),
                                .w_pr_gs_over      (      w_pr_gs_over_c1b0_gen[i]),
                                .w_pr_size_over    (    w_pr_size_over_c1b0_gen[i]),
                                .w_pr_0f           (           w_pr_0f_c1b0_gen[i]),
                                .w_pr_pos          (          w_pr_pos_c1b0_gen[i]),
                                .w_mux_sel         (         w_mux_sel_c1b0_gen[i]));
  end
endgenerate

mux_nbit_32x1 #3 u_mux_sel2(.a0  (w_mux_sel_c1b0_gen[0 ]),  
                           .a1  (w_mux_sel_c1b0_gen[1 ]),
                           .a2  (w_mux_sel_c1b0_gen[2 ]),
                           .a3  (w_mux_sel_c1b0_gen[3 ]),
                           .a4  (w_mux_sel_c1b0_gen[4 ]),
                           .a5  (w_mux_sel_c1b0_gen[5 ]),
                           .a6  (w_mux_sel_c1b0_gen[6 ]),
                           .a7  (w_mux_sel_c1b0_gen[7 ]),
                           .a8  (w_mux_sel_c1b0_gen[8 ]),
                           .a9  (w_mux_sel_c1b0_gen[9 ]),
                           .a10 (w_mux_sel_c1b0_gen[10]),
                           .a11 (w_mux_sel_c1b0_gen[11]),
                           .a12 (w_mux_sel_c1b0_gen[12]),
                           .a13 (w_mux_sel_c1b0_gen[13]),
                           .a14 (w_mux_sel_c1b0_gen[14]),
                           .a15 (w_mux_sel_c1b0_gen[15]),
                           .a16 (w_mux_sel_c1b0_gen[16]),
                           .a17 (w_mux_sel_c1b0_gen[17]),
                           .a18 (w_mux_sel_c1b0_gen[18]),
                           .a19 (w_mux_sel_c1b0_gen[19]),
                           .a20 (w_mux_sel_c1b0_gen[20]),
                           .a21 (w_mux_sel_c1b0_gen[21]),
                           .a22 (w_mux_sel_c1b0_gen[22]),
                           .a23 (w_mux_sel_c1b0_gen[23]),
                           .a24 (w_mux_sel_c1b0_gen[24]),
                           .a25 (w_mux_sel_c1b0_gen[25]),
                           .a26 (w_mux_sel_c1b0_gen[26]),
                           .a27 (w_mux_sel_c1b0_gen[27]),
                           .a28 (w_mux_sel_c1b0_gen[28]),
                           .a29 (w_mux_sel_c1b0_gen[29]),
                           .a30 (w_mux_sel_c1b0_gen[30]),
                           .a31 (w_mux_sel_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_mux_sel_c1b0));


mux_nbit_32x1 #4 u_pr_repn2(.a0  (w_pr_repne_c1b0_gen[0 ]),  
                           .a1  (w_pr_repne_c1b0_gen[1 ]),
                           .a2  (w_pr_repne_c1b0_gen[2 ]),
                           .a3  (w_pr_repne_c1b0_gen[3 ]),
                           .a4  (w_pr_repne_c1b0_gen[4 ]),
                           .a5  (w_pr_repne_c1b0_gen[5 ]),
                           .a6  (w_pr_repne_c1b0_gen[6 ]),
                           .a7  (w_pr_repne_c1b0_gen[7 ]),
                           .a8  (w_pr_repne_c1b0_gen[8 ]),
                           .a9  (w_pr_repne_c1b0_gen[9 ]),
                           .a10 (w_pr_repne_c1b0_gen[10]),
                           .a11 (w_pr_repne_c1b0_gen[11]),
                           .a12 (w_pr_repne_c1b0_gen[12]),
                           .a13 (w_pr_repne_c1b0_gen[13]),
                           .a14 (w_pr_repne_c1b0_gen[14]),
                           .a15 (w_pr_repne_c1b0_gen[15]),
                           .a16 (w_pr_repne_c1b0_gen[16]),
                           .a17 (w_pr_repne_c1b0_gen[17]),
                           .a18 (w_pr_repne_c1b0_gen[18]),
                           .a19 (w_pr_repne_c1b0_gen[19]),
                           .a20 (w_pr_repne_c1b0_gen[20]),
                           .a21 (w_pr_repne_c1b0_gen[21]),
                           .a22 (w_pr_repne_c1b0_gen[22]),
                           .a23 (w_pr_repne_c1b0_gen[23]),
                           .a24 (w_pr_repne_c1b0_gen[24]),
                           .a25 (w_pr_repne_c1b0_gen[25]),
                           .a26 (w_pr_repne_c1b0_gen[26]),
                           .a27 (w_pr_repne_c1b0_gen[27]),
                           .a28 (w_pr_repne_c1b0_gen[28]),
                           .a29 (w_pr_repne_c1b0_gen[29]),
                           .a30 (w_pr_repne_c1b0_gen[30]),
                           .a31 (w_pr_repne_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_repne_c1b0));


mux_nbit_32x1 #4 u_pr_cs2  (.a0  (w_pr_cs_over_c1b0_gen[0 ]),  
                           .a1  (w_pr_cs_over_c1b0_gen[1 ]),
                           .a2  (w_pr_cs_over_c1b0_gen[2 ]),
                           .a3  (w_pr_cs_over_c1b0_gen[3 ]),
                           .a4  (w_pr_cs_over_c1b0_gen[4 ]),
                           .a5  (w_pr_cs_over_c1b0_gen[5 ]),
                           .a6  (w_pr_cs_over_c1b0_gen[6 ]),
                           .a7  (w_pr_cs_over_c1b0_gen[7 ]),
                           .a8  (w_pr_cs_over_c1b0_gen[8 ]),
                           .a9  (w_pr_cs_over_c1b0_gen[9 ]),
                           .a10 (w_pr_cs_over_c1b0_gen[10]),
                           .a11 (w_pr_cs_over_c1b0_gen[11]),
                           .a12 (w_pr_cs_over_c1b0_gen[12]),
                           .a13 (w_pr_cs_over_c1b0_gen[13]),
                           .a14 (w_pr_cs_over_c1b0_gen[14]),
                           .a15 (w_pr_cs_over_c1b0_gen[15]),
                           .a16 (w_pr_cs_over_c1b0_gen[16]),
                           .a17 (w_pr_cs_over_c1b0_gen[17]),
                           .a18 (w_pr_cs_over_c1b0_gen[18]),
                           .a19 (w_pr_cs_over_c1b0_gen[19]),
                           .a20 (w_pr_cs_over_c1b0_gen[20]),
                           .a21 (w_pr_cs_over_c1b0_gen[21]),
                           .a22 (w_pr_cs_over_c1b0_gen[22]),
                           .a23 (w_pr_cs_over_c1b0_gen[23]),
                           .a24 (w_pr_cs_over_c1b0_gen[24]),
                           .a25 (w_pr_cs_over_c1b0_gen[25]),
                           .a26 (w_pr_cs_over_c1b0_gen[26]),
                           .a27 (w_pr_cs_over_c1b0_gen[27]),
                           .a28 (w_pr_cs_over_c1b0_gen[28]),
                           .a29 (w_pr_cs_over_c1b0_gen[29]),
                           .a30 (w_pr_cs_over_c1b0_gen[30]),
                           .a31 (w_pr_cs_over_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_cs_over_c1b0));

mux_nbit_32x1 #4 u_pr_ss2  (.a0  (w_pr_ss_over_c1b0_gen[0 ]),  
                           .a1  (w_pr_ss_over_c1b0_gen[1 ]),
                           .a2  (w_pr_ss_over_c1b0_gen[2 ]),
                           .a3  (w_pr_ss_over_c1b0_gen[3 ]),
                           .a4  (w_pr_ss_over_c1b0_gen[4 ]),
                           .a5  (w_pr_ss_over_c1b0_gen[5 ]),
                           .a6  (w_pr_ss_over_c1b0_gen[6 ]),
                           .a7  (w_pr_ss_over_c1b0_gen[7 ]),
                           .a8  (w_pr_ss_over_c1b0_gen[8 ]),
                           .a9  (w_pr_ss_over_c1b0_gen[9 ]),
                           .a10 (w_pr_ss_over_c1b0_gen[10]),
                           .a11 (w_pr_ss_over_c1b0_gen[11]),
                           .a12 (w_pr_ss_over_c1b0_gen[12]),
                           .a13 (w_pr_ss_over_c1b0_gen[13]),
                           .a14 (w_pr_ss_over_c1b0_gen[14]),
                           .a15 (w_pr_ss_over_c1b0_gen[15]),
                           .a16 (w_pr_ss_over_c1b0_gen[16]),
                           .a17 (w_pr_ss_over_c1b0_gen[17]),
                           .a18 (w_pr_ss_over_c1b0_gen[18]),
                           .a19 (w_pr_ss_over_c1b0_gen[19]),
                           .a20 (w_pr_ss_over_c1b0_gen[20]),
                           .a21 (w_pr_ss_over_c1b0_gen[21]),
                           .a22 (w_pr_ss_over_c1b0_gen[22]),
                           .a23 (w_pr_ss_over_c1b0_gen[23]),
                           .a24 (w_pr_ss_over_c1b0_gen[24]),
                           .a25 (w_pr_ss_over_c1b0_gen[25]),
                           .a26 (w_pr_ss_over_c1b0_gen[26]),
                           .a27 (w_pr_ss_over_c1b0_gen[27]),
                           .a28 (w_pr_ss_over_c1b0_gen[28]),
                           .a29 (w_pr_ss_over_c1b0_gen[29]),
                           .a30 (w_pr_ss_over_c1b0_gen[30]),
                           .a31 (w_pr_ss_over_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ss_over_c1b0));

mux_nbit_32x1 #4 u_pr_ds2  (.a0  (w_pr_ds_over_c1b0_gen[0 ]),  
                           .a1  (w_pr_ds_over_c1b0_gen[1 ]),
                           .a2  (w_pr_ds_over_c1b0_gen[2 ]),
                           .a3  (w_pr_ds_over_c1b0_gen[3 ]),
                           .a4  (w_pr_ds_over_c1b0_gen[4 ]),
                           .a5  (w_pr_ds_over_c1b0_gen[5 ]),
                           .a6  (w_pr_ds_over_c1b0_gen[6 ]),
                           .a7  (w_pr_ds_over_c1b0_gen[7 ]),
                           .a8  (w_pr_ds_over_c1b0_gen[8 ]),
                           .a9  (w_pr_ds_over_c1b0_gen[9 ]),
                           .a10 (w_pr_ds_over_c1b0_gen[10]),
                           .a11 (w_pr_ds_over_c1b0_gen[11]),
                           .a12 (w_pr_ds_over_c1b0_gen[12]),
                           .a13 (w_pr_ds_over_c1b0_gen[13]),
                           .a14 (w_pr_ds_over_c1b0_gen[14]),
                           .a15 (w_pr_ds_over_c1b0_gen[15]),
                           .a16 (w_pr_ds_over_c1b0_gen[16]),
                           .a17 (w_pr_ds_over_c1b0_gen[17]),
                           .a18 (w_pr_ds_over_c1b0_gen[18]),
                           .a19 (w_pr_ds_over_c1b0_gen[19]),
                           .a20 (w_pr_ds_over_c1b0_gen[20]),
                           .a21 (w_pr_ds_over_c1b0_gen[21]),
                           .a22 (w_pr_ds_over_c1b0_gen[22]),
                           .a23 (w_pr_ds_over_c1b0_gen[23]),
                           .a24 (w_pr_ds_over_c1b0_gen[24]),
                           .a25 (w_pr_ds_over_c1b0_gen[25]),
                           .a26 (w_pr_ds_over_c1b0_gen[26]),
                           .a27 (w_pr_ds_over_c1b0_gen[27]),
                           .a28 (w_pr_ds_over_c1b0_gen[28]),
                           .a29 (w_pr_ds_over_c1b0_gen[29]),
                           .a30 (w_pr_ds_over_c1b0_gen[30]),
                           .a31 (w_pr_ds_over_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ds_over_c1b0));

mux_nbit_32x1 #4 u_pr_es2  (.a0  (w_pr_es_over_c1b0_gen[0 ]),  
                           .a1  (w_pr_es_over_c1b0_gen[1 ]),
                           .a2  (w_pr_es_over_c1b0_gen[2 ]),
                           .a3  (w_pr_es_over_c1b0_gen[3 ]),
                           .a4  (w_pr_es_over_c1b0_gen[4 ]),
                           .a5  (w_pr_es_over_c1b0_gen[5 ]),
                           .a6  (w_pr_es_over_c1b0_gen[6 ]),
                           .a7  (w_pr_es_over_c1b0_gen[7 ]),
                           .a8  (w_pr_es_over_c1b0_gen[8 ]),
                           .a9  (w_pr_es_over_c1b0_gen[9 ]),
                           .a10 (w_pr_es_over_c1b0_gen[10]),
                           .a11 (w_pr_es_over_c1b0_gen[11]),
                           .a12 (w_pr_es_over_c1b0_gen[12]),
                           .a13 (w_pr_es_over_c1b0_gen[13]),
                           .a14 (w_pr_es_over_c1b0_gen[14]),
                           .a15 (w_pr_es_over_c1b0_gen[15]),
                           .a16 (w_pr_es_over_c1b0_gen[16]),
                           .a17 (w_pr_es_over_c1b0_gen[17]),
                           .a18 (w_pr_es_over_c1b0_gen[18]),
                           .a19 (w_pr_es_over_c1b0_gen[19]),
                           .a20 (w_pr_es_over_c1b0_gen[20]),
                           .a21 (w_pr_es_over_c1b0_gen[21]),
                           .a22 (w_pr_es_over_c1b0_gen[22]),
                           .a23 (w_pr_es_over_c1b0_gen[23]),
                           .a24 (w_pr_es_over_c1b0_gen[24]),
                           .a25 (w_pr_es_over_c1b0_gen[25]),
                           .a26 (w_pr_es_over_c1b0_gen[26]),
                           .a27 (w_pr_es_over_c1b0_gen[27]),
                           .a28 (w_pr_es_over_c1b0_gen[28]),
                           .a29 (w_pr_es_over_c1b0_gen[29]),
                           .a30 (w_pr_es_over_c1b0_gen[30]),
                           .a31 (w_pr_es_over_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_es_over_c1b0));

mux_nbit_32x1 #4 u_pr_fs2  (.a0  (w_pr_fs_over_c1b0_gen[0 ]),  
                           .a1  (w_pr_fs_over_c1b0_gen[1 ]),
                           .a2  (w_pr_fs_over_c1b0_gen[2 ]),
                           .a3  (w_pr_fs_over_c1b0_gen[3 ]),
                           .a4  (w_pr_fs_over_c1b0_gen[4 ]),
                           .a5  (w_pr_fs_over_c1b0_gen[5 ]),
                           .a6  (w_pr_fs_over_c1b0_gen[6 ]),
                           .a7  (w_pr_fs_over_c1b0_gen[7 ]),
                           .a8  (w_pr_fs_over_c1b0_gen[8 ]),
                           .a9  (w_pr_fs_over_c1b0_gen[9 ]),
                           .a10 (w_pr_fs_over_c1b0_gen[10]),
                           .a11 (w_pr_fs_over_c1b0_gen[11]),
                           .a12 (w_pr_fs_over_c1b0_gen[12]),
                           .a13 (w_pr_fs_over_c1b0_gen[13]),
                           .a14 (w_pr_fs_over_c1b0_gen[14]),
                           .a15 (w_pr_fs_over_c1b0_gen[15]),
                           .a16 (w_pr_fs_over_c1b0_gen[16]),
                           .a17 (w_pr_fs_over_c1b0_gen[17]),
                           .a18 (w_pr_fs_over_c1b0_gen[18]),
                           .a19 (w_pr_fs_over_c1b0_gen[19]),
                           .a20 (w_pr_fs_over_c1b0_gen[20]),
                           .a21 (w_pr_fs_over_c1b0_gen[21]),
                           .a22 (w_pr_fs_over_c1b0_gen[22]),
                           .a23 (w_pr_fs_over_c1b0_gen[23]),
                           .a24 (w_pr_fs_over_c1b0_gen[24]),
                           .a25 (w_pr_fs_over_c1b0_gen[25]),
                           .a26 (w_pr_fs_over_c1b0_gen[26]),
                           .a27 (w_pr_fs_over_c1b0_gen[27]),
                           .a28 (w_pr_fs_over_c1b0_gen[28]),
                           .a29 (w_pr_fs_over_c1b0_gen[29]),
                           .a30 (w_pr_fs_over_c1b0_gen[30]),
                           .a31 (w_pr_fs_over_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_fs_over_c1b0));

mux_nbit_32x1 #4 u_pr_gs2  (.a0  (w_pr_gs_over_c1b0_gen[0 ]),  
                           .a1  (w_pr_gs_over_c1b0_gen[1 ]),
                           .a2  (w_pr_gs_over_c1b0_gen[2 ]),
                           .a3  (w_pr_gs_over_c1b0_gen[3 ]),
                           .a4  (w_pr_gs_over_c1b0_gen[4 ]),
                           .a5  (w_pr_gs_over_c1b0_gen[5 ]),
                           .a6  (w_pr_gs_over_c1b0_gen[6 ]),
                           .a7  (w_pr_gs_over_c1b0_gen[7 ]),
                           .a8  (w_pr_gs_over_c1b0_gen[8 ]),
                           .a9  (w_pr_gs_over_c1b0_gen[9 ]),
                           .a10 (w_pr_gs_over_c1b0_gen[10]),
                           .a11 (w_pr_gs_over_c1b0_gen[11]),
                           .a12 (w_pr_gs_over_c1b0_gen[12]),
                           .a13 (w_pr_gs_over_c1b0_gen[13]),
                           .a14 (w_pr_gs_over_c1b0_gen[14]),
                           .a15 (w_pr_gs_over_c1b0_gen[15]),
                           .a16 (w_pr_gs_over_c1b0_gen[16]),
                           .a17 (w_pr_gs_over_c1b0_gen[17]),
                           .a18 (w_pr_gs_over_c1b0_gen[18]),
                           .a19 (w_pr_gs_over_c1b0_gen[19]),
                           .a20 (w_pr_gs_over_c1b0_gen[20]),
                           .a21 (w_pr_gs_over_c1b0_gen[21]),
                           .a22 (w_pr_gs_over_c1b0_gen[22]),
                           .a23 (w_pr_gs_over_c1b0_gen[23]),
                           .a24 (w_pr_gs_over_c1b0_gen[24]),
                           .a25 (w_pr_gs_over_c1b0_gen[25]),
                           .a26 (w_pr_gs_over_c1b0_gen[26]),
                           .a27 (w_pr_gs_over_c1b0_gen[27]),
                           .a28 (w_pr_gs_over_c1b0_gen[28]),
                           .a29 (w_pr_gs_over_c1b0_gen[29]),
                           .a30 (w_pr_gs_over_c1b0_gen[30]),
                           .a31 (w_pr_gs_over_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_gs_over_c1b0));

mux_nbit_32x1 #4 u_pr_size2(.a0  (w_pr_size_over_c1b0_gen[0 ]),  
                           .a1  (w_pr_size_over_c1b0_gen[1 ]),
                           .a2  (w_pr_size_over_c1b0_gen[2 ]),
                           .a3  (w_pr_size_over_c1b0_gen[3 ]),
                           .a4  (w_pr_size_over_c1b0_gen[4 ]),
                           .a5  (w_pr_size_over_c1b0_gen[5 ]),
                           .a6  (w_pr_size_over_c1b0_gen[6 ]),
                           .a7  (w_pr_size_over_c1b0_gen[7 ]),
                           .a8  (w_pr_size_over_c1b0_gen[8 ]),
                           .a9  (w_pr_size_over_c1b0_gen[9 ]),
                           .a10 (w_pr_size_over_c1b0_gen[10]),
                           .a11 (w_pr_size_over_c1b0_gen[11]),
                           .a12 (w_pr_size_over_c1b0_gen[12]),
                           .a13 (w_pr_size_over_c1b0_gen[13]),
                           .a14 (w_pr_size_over_c1b0_gen[14]),
                           .a15 (w_pr_size_over_c1b0_gen[15]),
                           .a16 (w_pr_size_over_c1b0_gen[16]),
                           .a17 (w_pr_size_over_c1b0_gen[17]),
                           .a18 (w_pr_size_over_c1b0_gen[18]),
                           .a19 (w_pr_size_over_c1b0_gen[19]),
                           .a20 (w_pr_size_over_c1b0_gen[20]),
                           .a21 (w_pr_size_over_c1b0_gen[21]),
                           .a22 (w_pr_size_over_c1b0_gen[22]),
                           .a23 (w_pr_size_over_c1b0_gen[23]),
                           .a24 (w_pr_size_over_c1b0_gen[24]),
                           .a25 (w_pr_size_over_c1b0_gen[25]),
                           .a26 (w_pr_size_over_c1b0_gen[26]),
                           .a27 (w_pr_size_over_c1b0_gen[27]),
                           .a28 (w_pr_size_over_c1b0_gen[28]),
                           .a29 (w_pr_size_over_c1b0_gen[29]),
                           .a30 (w_pr_size_over_c1b0_gen[30]),
                           .a31 (w_pr_size_over_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_size_over_c1b0));

mux_nbit_32x1 #4 u_pr_0f2  (.a0  (w_pr_0f_c1b0_gen[0 ]),  
                           .a1  (w_pr_0f_c1b0_gen[1 ]),
                           .a2  (w_pr_0f_c1b0_gen[2 ]),
                           .a3  (w_pr_0f_c1b0_gen[3 ]),
                           .a4  (w_pr_0f_c1b0_gen[4 ]),
                           .a5  (w_pr_0f_c1b0_gen[5 ]),
                           .a6  (w_pr_0f_c1b0_gen[6 ]),
                           .a7  (w_pr_0f_c1b0_gen[7 ]),
                           .a8  (w_pr_0f_c1b0_gen[8 ]),
                           .a9  (w_pr_0f_c1b0_gen[9 ]),
                           .a10 (w_pr_0f_c1b0_gen[10]),
                           .a11 (w_pr_0f_c1b0_gen[11]),
                           .a12 (w_pr_0f_c1b0_gen[12]),
                           .a13 (w_pr_0f_c1b0_gen[13]),
                           .a14 (w_pr_0f_c1b0_gen[14]),
                           .a15 (w_pr_0f_c1b0_gen[15]),
                           .a16 (w_pr_0f_c1b0_gen[16]),
                           .a17 (w_pr_0f_c1b0_gen[17]),
                           .a18 (w_pr_0f_c1b0_gen[18]),
                           .a19 (w_pr_0f_c1b0_gen[19]),
                           .a20 (w_pr_0f_c1b0_gen[20]),
                           .a21 (w_pr_0f_c1b0_gen[21]),
                           .a22 (w_pr_0f_c1b0_gen[22]),
                           .a23 (w_pr_0f_c1b0_gen[23]),
                           .a24 (w_pr_0f_c1b0_gen[24]),
                           .a25 (w_pr_0f_c1b0_gen[25]),
                           .a26 (w_pr_0f_c1b0_gen[26]),
                           .a27 (w_pr_0f_c1b0_gen[27]),
                           .a28 (w_pr_0f_c1b0_gen[28]),
                           .a29 (w_pr_0f_c1b0_gen[29]),
                           .a30 (w_pr_0f_c1b0_gen[30]),
                           .a31 (w_pr_0f_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_0f_c1b0));

mux_nbit_32x1 #4 u_pr_pos2  (.a0  (w_pr_pos_c1b0_gen[0 ]),  
                           .a1  (w_pr_pos_c1b0_gen[1 ]),
                           .a2  (w_pr_pos_c1b0_gen[2 ]),
                           .a3  (w_pr_pos_c1b0_gen[3 ]),
                           .a4  (w_pr_pos_c1b0_gen[4 ]),
                           .a5  (w_pr_pos_c1b0_gen[5 ]),
                           .a6  (w_pr_pos_c1b0_gen[6 ]),
                           .a7  (w_pr_pos_c1b0_gen[7 ]),
                           .a8  (w_pr_pos_c1b0_gen[8 ]),
                           .a9  (w_pr_pos_c1b0_gen[9 ]),
                           .a10 (w_pr_pos_c1b0_gen[10]),
                           .a11 (w_pr_pos_c1b0_gen[11]),
                           .a12 (w_pr_pos_c1b0_gen[12]),
                           .a13 (w_pr_pos_c1b0_gen[13]),
                           .a14 (w_pr_pos_c1b0_gen[14]),
                           .a15 (w_pr_pos_c1b0_gen[15]),
                           .a16 (w_pr_pos_c1b0_gen[16]),
                           .a17 (w_pr_pos_c1b0_gen[17]),
                           .a18 (w_pr_pos_c1b0_gen[18]),
                           .a19 (w_pr_pos_c1b0_gen[19]),
                           .a20 (w_pr_pos_c1b0_gen[20]),
                           .a21 (w_pr_pos_c1b0_gen[21]),
                           .a22 (w_pr_pos_c1b0_gen[22]),
                           .a23 (w_pr_pos_c1b0_gen[23]),
                           .a24 (w_pr_pos_c1b0_gen[24]),
                           .a25 (w_pr_pos_c1b0_gen[25]),
                           .a26 (w_pr_pos_c1b0_gen[26]),
                           .a27 (w_pr_pos_c1b0_gen[27]),
                           .a28 (w_pr_pos_c1b0_gen[28]),
                           .a29 (w_pr_pos_c1b0_gen[29]),
                           .a30 (w_pr_pos_c1b0_gen[30]),
                           .a31 (w_pr_pos_c1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_pos_c1b0));
//b1c0
generate
  for (i=0; i<32; i=i+1) begin : fetch_dec3
fetch_to_decode u_fetch_decode3 (.de_lower_16bytes  (        b1c0[((i*8)+31):i*8]), 
                                .w_pr_repne        (        w_pr_repne_b1c0_gen[i]),
                                .w_pr_cs_over      (      w_pr_cs_over_b1c0_gen[i]),
                                .w_pr_ss_over      (      w_pr_ss_over_b1c0_gen[i]),
                                .w_pr_ds_over      (      w_pr_ds_over_b1c0_gen[i]),
                                .w_pr_es_over      (      w_pr_es_over_b1c0_gen[i]),
                                .w_pr_fs_over      (      w_pr_fs_over_b1c0_gen[i]),
                                .w_pr_gs_over      (      w_pr_gs_over_b1c0_gen[i]),
                                .w_pr_size_over    (    w_pr_size_over_b1c0_gen[i]),
                                .w_pr_0f           (           w_pr_0f_b1c0_gen[i]),
                                .w_pr_pos          (          w_pr_pos_b1c0_gen[i]),
                                .w_mux_sel         (         w_mux_sel_b1c0_gen[i]));
  end
endgenerate

mux_nbit_32x1 #3 u_mux_sel3(.a0  (w_mux_sel_b1c0_gen[0 ]),  
                           .a1  (w_mux_sel_b1c0_gen[1 ]),
                           .a2  (w_mux_sel_b1c0_gen[2 ]),
                           .a3  (w_mux_sel_b1c0_gen[3 ]),
                           .a4  (w_mux_sel_b1c0_gen[4 ]),
                           .a5  (w_mux_sel_b1c0_gen[5 ]),
                           .a6  (w_mux_sel_b1c0_gen[6 ]),
                           .a7  (w_mux_sel_b1c0_gen[7 ]),
                           .a8  (w_mux_sel_b1c0_gen[8 ]),
                           .a9  (w_mux_sel_b1c0_gen[9 ]),
                           .a10 (w_mux_sel_b1c0_gen[10]),
                           .a11 (w_mux_sel_b1c0_gen[11]),
                           .a12 (w_mux_sel_b1c0_gen[12]),
                           .a13 (w_mux_sel_b1c0_gen[13]),
                           .a14 (w_mux_sel_b1c0_gen[14]),
                           .a15 (w_mux_sel_b1c0_gen[15]),
                           .a16 (w_mux_sel_b1c0_gen[16]),
                           .a17 (w_mux_sel_b1c0_gen[17]),
                           .a18 (w_mux_sel_b1c0_gen[18]),
                           .a19 (w_mux_sel_b1c0_gen[19]),
                           .a20 (w_mux_sel_b1c0_gen[20]),
                           .a21 (w_mux_sel_b1c0_gen[21]),
                           .a22 (w_mux_sel_b1c0_gen[22]),
                           .a23 (w_mux_sel_b1c0_gen[23]),
                           .a24 (w_mux_sel_b1c0_gen[24]),
                           .a25 (w_mux_sel_b1c0_gen[25]),
                           .a26 (w_mux_sel_b1c0_gen[26]),
                           .a27 (w_mux_sel_b1c0_gen[27]),
                           .a28 (w_mux_sel_b1c0_gen[28]),
                           .a29 (w_mux_sel_b1c0_gen[29]),
                           .a30 (w_mux_sel_b1c0_gen[30]),
                           .a31 (w_mux_sel_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_mux_sel_b1c0));


mux_nbit_32x1 #4 u_pr_repn3(.a0  (w_pr_repne_b1c0_gen[0 ]),  
                           .a1  (w_pr_repne_b1c0_gen[1 ]),
                           .a2  (w_pr_repne_b1c0_gen[2 ]),
                           .a3  (w_pr_repne_b1c0_gen[3 ]),
                           .a4  (w_pr_repne_b1c0_gen[4 ]),
                           .a5  (w_pr_repne_b1c0_gen[5 ]),
                           .a6  (w_pr_repne_b1c0_gen[6 ]),
                           .a7  (w_pr_repne_b1c0_gen[7 ]),
                           .a8  (w_pr_repne_b1c0_gen[8 ]),
                           .a9  (w_pr_repne_b1c0_gen[9 ]),
                           .a10 (w_pr_repne_b1c0_gen[10]),
                           .a11 (w_pr_repne_b1c0_gen[11]),
                           .a12 (w_pr_repne_b1c0_gen[12]),
                           .a13 (w_pr_repne_b1c0_gen[13]),
                           .a14 (w_pr_repne_b1c0_gen[14]),
                           .a15 (w_pr_repne_b1c0_gen[15]),
                           .a16 (w_pr_repne_b1c0_gen[16]),
                           .a17 (w_pr_repne_b1c0_gen[17]),
                           .a18 (w_pr_repne_b1c0_gen[18]),
                           .a19 (w_pr_repne_b1c0_gen[19]),
                           .a20 (w_pr_repne_b1c0_gen[20]),
                           .a21 (w_pr_repne_b1c0_gen[21]),
                           .a22 (w_pr_repne_b1c0_gen[22]),
                           .a23 (w_pr_repne_b1c0_gen[23]),
                           .a24 (w_pr_repne_b1c0_gen[24]),
                           .a25 (w_pr_repne_b1c0_gen[25]),
                           .a26 (w_pr_repne_b1c0_gen[26]),
                           .a27 (w_pr_repne_b1c0_gen[27]),
                           .a28 (w_pr_repne_b1c0_gen[28]),
                           .a29 (w_pr_repne_b1c0_gen[29]),
                           .a30 (w_pr_repne_b1c0_gen[30]),
                           .a31 (w_pr_repne_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_repne_b1c0));


mux_nbit_32x1 #4 u_pr_cs3  (.a0  (w_pr_cs_over_b1c0_gen[0 ]),  
                           .a1  (w_pr_cs_over_b1c0_gen[1 ]),
                           .a2  (w_pr_cs_over_b1c0_gen[2 ]),
                           .a3  (w_pr_cs_over_b1c0_gen[3 ]),
                           .a4  (w_pr_cs_over_b1c0_gen[4 ]),
                           .a5  (w_pr_cs_over_b1c0_gen[5 ]),
                           .a6  (w_pr_cs_over_b1c0_gen[6 ]),
                           .a7  (w_pr_cs_over_b1c0_gen[7 ]),
                           .a8  (w_pr_cs_over_b1c0_gen[8 ]),
                           .a9  (w_pr_cs_over_b1c0_gen[9 ]),
                           .a10 (w_pr_cs_over_b1c0_gen[10]),
                           .a11 (w_pr_cs_over_b1c0_gen[11]),
                           .a12 (w_pr_cs_over_b1c0_gen[12]),
                           .a13 (w_pr_cs_over_b1c0_gen[13]),
                           .a14 (w_pr_cs_over_b1c0_gen[14]),
                           .a15 (w_pr_cs_over_b1c0_gen[15]),
                           .a16 (w_pr_cs_over_b1c0_gen[16]),
                           .a17 (w_pr_cs_over_b1c0_gen[17]),
                           .a18 (w_pr_cs_over_b1c0_gen[18]),
                           .a19 (w_pr_cs_over_b1c0_gen[19]),
                           .a20 (w_pr_cs_over_b1c0_gen[20]),
                           .a21 (w_pr_cs_over_b1c0_gen[21]),
                           .a22 (w_pr_cs_over_b1c0_gen[22]),
                           .a23 (w_pr_cs_over_b1c0_gen[23]),
                           .a24 (w_pr_cs_over_b1c0_gen[24]),
                           .a25 (w_pr_cs_over_b1c0_gen[25]),
                           .a26 (w_pr_cs_over_b1c0_gen[26]),
                           .a27 (w_pr_cs_over_b1c0_gen[27]),
                           .a28 (w_pr_cs_over_b1c0_gen[28]),
                           .a29 (w_pr_cs_over_b1c0_gen[29]),
                           .a30 (w_pr_cs_over_b1c0_gen[30]),
                           .a31 (w_pr_cs_over_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_cs_over_b1c0));

mux_nbit_32x1 #4 u_pr_ss3  (.a0  (w_pr_ss_over_b1c0_gen[0 ]),  
                           .a1  (w_pr_ss_over_b1c0_gen[1 ]),
                           .a2  (w_pr_ss_over_b1c0_gen[2 ]),
                           .a3  (w_pr_ss_over_b1c0_gen[3 ]),
                           .a4  (w_pr_ss_over_b1c0_gen[4 ]),
                           .a5  (w_pr_ss_over_b1c0_gen[5 ]),
                           .a6  (w_pr_ss_over_b1c0_gen[6 ]),
                           .a7  (w_pr_ss_over_b1c0_gen[7 ]),
                           .a8  (w_pr_ss_over_b1c0_gen[8 ]),
                           .a9  (w_pr_ss_over_b1c0_gen[9 ]),
                           .a10 (w_pr_ss_over_b1c0_gen[10]),
                           .a11 (w_pr_ss_over_b1c0_gen[11]),
                           .a12 (w_pr_ss_over_b1c0_gen[12]),
                           .a13 (w_pr_ss_over_b1c0_gen[13]),
                           .a14 (w_pr_ss_over_b1c0_gen[14]),
                           .a15 (w_pr_ss_over_b1c0_gen[15]),
                           .a16 (w_pr_ss_over_b1c0_gen[16]),
                           .a17 (w_pr_ss_over_b1c0_gen[17]),
                           .a18 (w_pr_ss_over_b1c0_gen[18]),
                           .a19 (w_pr_ss_over_b1c0_gen[19]),
                           .a20 (w_pr_ss_over_b1c0_gen[20]),
                           .a21 (w_pr_ss_over_b1c0_gen[21]),
                           .a22 (w_pr_ss_over_b1c0_gen[22]),
                           .a23 (w_pr_ss_over_b1c0_gen[23]),
                           .a24 (w_pr_ss_over_b1c0_gen[24]),
                           .a25 (w_pr_ss_over_b1c0_gen[25]),
                           .a26 (w_pr_ss_over_b1c0_gen[26]),
                           .a27 (w_pr_ss_over_b1c0_gen[27]),
                           .a28 (w_pr_ss_over_b1c0_gen[28]),
                           .a29 (w_pr_ss_over_b1c0_gen[29]),
                           .a30 (w_pr_ss_over_b1c0_gen[30]),
                           .a31 (w_pr_ss_over_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ss_over_b1c0));

mux_nbit_32x1 #4 u_pr_ds3  (.a0  (w_pr_ds_over_b1c0_gen[0 ]),  
                           .a1  (w_pr_ds_over_b1c0_gen[1 ]),
                           .a2  (w_pr_ds_over_b1c0_gen[2 ]),
                           .a3  (w_pr_ds_over_b1c0_gen[3 ]),
                           .a4  (w_pr_ds_over_b1c0_gen[4 ]),
                           .a5  (w_pr_ds_over_b1c0_gen[5 ]),
                           .a6  (w_pr_ds_over_b1c0_gen[6 ]),
                           .a7  (w_pr_ds_over_b1c0_gen[7 ]),
                           .a8  (w_pr_ds_over_b1c0_gen[8 ]),
                           .a9  (w_pr_ds_over_b1c0_gen[9 ]),
                           .a10 (w_pr_ds_over_b1c0_gen[10]),
                           .a11 (w_pr_ds_over_b1c0_gen[11]),
                           .a12 (w_pr_ds_over_b1c0_gen[12]),
                           .a13 (w_pr_ds_over_b1c0_gen[13]),
                           .a14 (w_pr_ds_over_b1c0_gen[14]),
                           .a15 (w_pr_ds_over_b1c0_gen[15]),
                           .a16 (w_pr_ds_over_b1c0_gen[16]),
                           .a17 (w_pr_ds_over_b1c0_gen[17]),
                           .a18 (w_pr_ds_over_b1c0_gen[18]),
                           .a19 (w_pr_ds_over_b1c0_gen[19]),
                           .a20 (w_pr_ds_over_b1c0_gen[20]),
                           .a21 (w_pr_ds_over_b1c0_gen[21]),
                           .a22 (w_pr_ds_over_b1c0_gen[22]),
                           .a23 (w_pr_ds_over_b1c0_gen[23]),
                           .a24 (w_pr_ds_over_b1c0_gen[24]),
                           .a25 (w_pr_ds_over_b1c0_gen[25]),
                           .a26 (w_pr_ds_over_b1c0_gen[26]),
                           .a27 (w_pr_ds_over_b1c0_gen[27]),
                           .a28 (w_pr_ds_over_b1c0_gen[28]),
                           .a29 (w_pr_ds_over_b1c0_gen[29]),
                           .a30 (w_pr_ds_over_b1c0_gen[30]),
                           .a31 (w_pr_ds_over_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ds_over_b1c0));

mux_nbit_32x1 #4 u_pr_es3  (.a0  (w_pr_es_over_b1c0_gen[0 ]),  
                           .a1  (w_pr_es_over_b1c0_gen[1 ]),
                           .a2  (w_pr_es_over_b1c0_gen[2 ]),
                           .a3  (w_pr_es_over_b1c0_gen[3 ]),
                           .a4  (w_pr_es_over_b1c0_gen[4 ]),
                           .a5  (w_pr_es_over_b1c0_gen[5 ]),
                           .a6  (w_pr_es_over_b1c0_gen[6 ]),
                           .a7  (w_pr_es_over_b1c0_gen[7 ]),
                           .a8  (w_pr_es_over_b1c0_gen[8 ]),
                           .a9  (w_pr_es_over_b1c0_gen[9 ]),
                           .a10 (w_pr_es_over_b1c0_gen[10]),
                           .a11 (w_pr_es_over_b1c0_gen[11]),
                           .a12 (w_pr_es_over_b1c0_gen[12]),
                           .a13 (w_pr_es_over_b1c0_gen[13]),
                           .a14 (w_pr_es_over_b1c0_gen[14]),
                           .a15 (w_pr_es_over_b1c0_gen[15]),
                           .a16 (w_pr_es_over_b1c0_gen[16]),
                           .a17 (w_pr_es_over_b1c0_gen[17]),
                           .a18 (w_pr_es_over_b1c0_gen[18]),
                           .a19 (w_pr_es_over_b1c0_gen[19]),
                           .a20 (w_pr_es_over_b1c0_gen[20]),
                           .a21 (w_pr_es_over_b1c0_gen[21]),
                           .a22 (w_pr_es_over_b1c0_gen[22]),
                           .a23 (w_pr_es_over_b1c0_gen[23]),
                           .a24 (w_pr_es_over_b1c0_gen[24]),
                           .a25 (w_pr_es_over_b1c0_gen[25]),
                           .a26 (w_pr_es_over_b1c0_gen[26]),
                           .a27 (w_pr_es_over_b1c0_gen[27]),
                           .a28 (w_pr_es_over_b1c0_gen[28]),
                           .a29 (w_pr_es_over_b1c0_gen[29]),
                           .a30 (w_pr_es_over_b1c0_gen[30]),
                           .a31 (w_pr_es_over_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_es_over_b1c0));

mux_nbit_32x1 #4 u_pr_fs3  (.a0  (w_pr_fs_over_b1c0_gen[0 ]),  
                           .a1  (w_pr_fs_over_b1c0_gen[1 ]),
                           .a2  (w_pr_fs_over_b1c0_gen[2 ]),
                           .a3  (w_pr_fs_over_b1c0_gen[3 ]),
                           .a4  (w_pr_fs_over_b1c0_gen[4 ]),
                           .a5  (w_pr_fs_over_b1c0_gen[5 ]),
                           .a6  (w_pr_fs_over_b1c0_gen[6 ]),
                           .a7  (w_pr_fs_over_b1c0_gen[7 ]),
                           .a8  (w_pr_fs_over_b1c0_gen[8 ]),
                           .a9  (w_pr_fs_over_b1c0_gen[9 ]),
                           .a10 (w_pr_fs_over_b1c0_gen[10]),
                           .a11 (w_pr_fs_over_b1c0_gen[11]),
                           .a12 (w_pr_fs_over_b1c0_gen[12]),
                           .a13 (w_pr_fs_over_b1c0_gen[13]),
                           .a14 (w_pr_fs_over_b1c0_gen[14]),
                           .a15 (w_pr_fs_over_b1c0_gen[15]),
                           .a16 (w_pr_fs_over_b1c0_gen[16]),
                           .a17 (w_pr_fs_over_b1c0_gen[17]),
                           .a18 (w_pr_fs_over_b1c0_gen[18]),
                           .a19 (w_pr_fs_over_b1c0_gen[19]),
                           .a20 (w_pr_fs_over_b1c0_gen[20]),
                           .a21 (w_pr_fs_over_b1c0_gen[21]),
                           .a22 (w_pr_fs_over_b1c0_gen[22]),
                           .a23 (w_pr_fs_over_b1c0_gen[23]),
                           .a24 (w_pr_fs_over_b1c0_gen[24]),
                           .a25 (w_pr_fs_over_b1c0_gen[25]),
                           .a26 (w_pr_fs_over_b1c0_gen[26]),
                           .a27 (w_pr_fs_over_b1c0_gen[27]),
                           .a28 (w_pr_fs_over_b1c0_gen[28]),
                           .a29 (w_pr_fs_over_b1c0_gen[29]),
                           .a30 (w_pr_fs_over_b1c0_gen[30]),
                           .a31 (w_pr_fs_over_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_fs_over_b1c0));

mux_nbit_32x1 #4 u_pr_gs3  (.a0  (w_pr_gs_over_b1c0_gen[0 ]),  
                           .a1  (w_pr_gs_over_b1c0_gen[1 ]),
                           .a2  (w_pr_gs_over_b1c0_gen[2 ]),
                           .a3  (w_pr_gs_over_b1c0_gen[3 ]),
                           .a4  (w_pr_gs_over_b1c0_gen[4 ]),
                           .a5  (w_pr_gs_over_b1c0_gen[5 ]),
                           .a6  (w_pr_gs_over_b1c0_gen[6 ]),
                           .a7  (w_pr_gs_over_b1c0_gen[7 ]),
                           .a8  (w_pr_gs_over_b1c0_gen[8 ]),
                           .a9  (w_pr_gs_over_b1c0_gen[9 ]),
                           .a10 (w_pr_gs_over_b1c0_gen[10]),
                           .a11 (w_pr_gs_over_b1c0_gen[11]),
                           .a12 (w_pr_gs_over_b1c0_gen[12]),
                           .a13 (w_pr_gs_over_b1c0_gen[13]),
                           .a14 (w_pr_gs_over_b1c0_gen[14]),
                           .a15 (w_pr_gs_over_b1c0_gen[15]),
                           .a16 (w_pr_gs_over_b1c0_gen[16]),
                           .a17 (w_pr_gs_over_b1c0_gen[17]),
                           .a18 (w_pr_gs_over_b1c0_gen[18]),
                           .a19 (w_pr_gs_over_b1c0_gen[19]),
                           .a20 (w_pr_gs_over_b1c0_gen[20]),
                           .a21 (w_pr_gs_over_b1c0_gen[21]),
                           .a22 (w_pr_gs_over_b1c0_gen[22]),
                           .a23 (w_pr_gs_over_b1c0_gen[23]),
                           .a24 (w_pr_gs_over_b1c0_gen[24]),
                           .a25 (w_pr_gs_over_b1c0_gen[25]),
                           .a26 (w_pr_gs_over_b1c0_gen[26]),
                           .a27 (w_pr_gs_over_b1c0_gen[27]),
                           .a28 (w_pr_gs_over_b1c0_gen[28]),
                           .a29 (w_pr_gs_over_b1c0_gen[29]),
                           .a30 (w_pr_gs_over_b1c0_gen[30]),
                           .a31 (w_pr_gs_over_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_gs_over_b1c0));

mux_nbit_32x1 #4 u_pr_size3(.a0  (w_pr_size_over_b1c0_gen[0 ]),  
                           .a1  (w_pr_size_over_b1c0_gen[1 ]),
                           .a2  (w_pr_size_over_b1c0_gen[2 ]),
                           .a3  (w_pr_size_over_b1c0_gen[3 ]),
                           .a4  (w_pr_size_over_b1c0_gen[4 ]),
                           .a5  (w_pr_size_over_b1c0_gen[5 ]),
                           .a6  (w_pr_size_over_b1c0_gen[6 ]),
                           .a7  (w_pr_size_over_b1c0_gen[7 ]),
                           .a8  (w_pr_size_over_b1c0_gen[8 ]),
                           .a9  (w_pr_size_over_b1c0_gen[9 ]),
                           .a10 (w_pr_size_over_b1c0_gen[10]),
                           .a11 (w_pr_size_over_b1c0_gen[11]),
                           .a12 (w_pr_size_over_b1c0_gen[12]),
                           .a13 (w_pr_size_over_b1c0_gen[13]),
                           .a14 (w_pr_size_over_b1c0_gen[14]),
                           .a15 (w_pr_size_over_b1c0_gen[15]),
                           .a16 (w_pr_size_over_b1c0_gen[16]),
                           .a17 (w_pr_size_over_b1c0_gen[17]),
                           .a18 (w_pr_size_over_b1c0_gen[18]),
                           .a19 (w_pr_size_over_b1c0_gen[19]),
                           .a20 (w_pr_size_over_b1c0_gen[20]),
                           .a21 (w_pr_size_over_b1c0_gen[21]),
                           .a22 (w_pr_size_over_b1c0_gen[22]),
                           .a23 (w_pr_size_over_b1c0_gen[23]),
                           .a24 (w_pr_size_over_b1c0_gen[24]),
                           .a25 (w_pr_size_over_b1c0_gen[25]),
                           .a26 (w_pr_size_over_b1c0_gen[26]),
                           .a27 (w_pr_size_over_b1c0_gen[27]),
                           .a28 (w_pr_size_over_b1c0_gen[28]),
                           .a29 (w_pr_size_over_b1c0_gen[29]),
                           .a30 (w_pr_size_over_b1c0_gen[30]),
                           .a31 (w_pr_size_over_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_size_over_b1c0));

mux_nbit_32x1 #4 u_pr_0f3  (.a0  (w_pr_0f_b1c0_gen[0 ]),  
                           .a1  (w_pr_0f_b1c0_gen[1 ]),
                           .a2  (w_pr_0f_b1c0_gen[2 ]),
                           .a3  (w_pr_0f_b1c0_gen[3 ]),
                           .a4  (w_pr_0f_b1c0_gen[4 ]),
                           .a5  (w_pr_0f_b1c0_gen[5 ]),
                           .a6  (w_pr_0f_b1c0_gen[6 ]),
                           .a7  (w_pr_0f_b1c0_gen[7 ]),
                           .a8  (w_pr_0f_b1c0_gen[8 ]),
                           .a9  (w_pr_0f_b1c0_gen[9 ]),
                           .a10 (w_pr_0f_b1c0_gen[10]),
                           .a11 (w_pr_0f_b1c0_gen[11]),
                           .a12 (w_pr_0f_b1c0_gen[12]),
                           .a13 (w_pr_0f_b1c0_gen[13]),
                           .a14 (w_pr_0f_b1c0_gen[14]),
                           .a15 (w_pr_0f_b1c0_gen[15]),
                           .a16 (w_pr_0f_b1c0_gen[16]),
                           .a17 (w_pr_0f_b1c0_gen[17]),
                           .a18 (w_pr_0f_b1c0_gen[18]),
                           .a19 (w_pr_0f_b1c0_gen[19]),
                           .a20 (w_pr_0f_b1c0_gen[20]),
                           .a21 (w_pr_0f_b1c0_gen[21]),
                           .a22 (w_pr_0f_b1c0_gen[22]),
                           .a23 (w_pr_0f_b1c0_gen[23]),
                           .a24 (w_pr_0f_b1c0_gen[24]),
                           .a25 (w_pr_0f_b1c0_gen[25]),
                           .a26 (w_pr_0f_b1c0_gen[26]),
                           .a27 (w_pr_0f_b1c0_gen[27]),
                           .a28 (w_pr_0f_b1c0_gen[28]),
                           .a29 (w_pr_0f_b1c0_gen[29]),
                           .a30 (w_pr_0f_b1c0_gen[30]),
                           .a31 (w_pr_0f_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_0f_b1c0));

mux_nbit_32x1 #4 u_pr_pos3  (.a0  (w_pr_pos_b1c0_gen[0 ]),  
                           .a1  (w_pr_pos_b1c0_gen[1 ]),
                           .a2  (w_pr_pos_b1c0_gen[2 ]),
                           .a3  (w_pr_pos_b1c0_gen[3 ]),
                           .a4  (w_pr_pos_b1c0_gen[4 ]),
                           .a5  (w_pr_pos_b1c0_gen[5 ]),
                           .a6  (w_pr_pos_b1c0_gen[6 ]),
                           .a7  (w_pr_pos_b1c0_gen[7 ]),
                           .a8  (w_pr_pos_b1c0_gen[8 ]),
                           .a9  (w_pr_pos_b1c0_gen[9 ]),
                           .a10 (w_pr_pos_b1c0_gen[10]),
                           .a11 (w_pr_pos_b1c0_gen[11]),
                           .a12 (w_pr_pos_b1c0_gen[12]),
                           .a13 (w_pr_pos_b1c0_gen[13]),
                           .a14 (w_pr_pos_b1c0_gen[14]),
                           .a15 (w_pr_pos_b1c0_gen[15]),
                           .a16 (w_pr_pos_b1c0_gen[16]),
                           .a17 (w_pr_pos_b1c0_gen[17]),
                           .a18 (w_pr_pos_b1c0_gen[18]),
                           .a19 (w_pr_pos_b1c0_gen[19]),
                           .a20 (w_pr_pos_b1c0_gen[20]),
                           .a21 (w_pr_pos_b1c0_gen[21]),
                           .a22 (w_pr_pos_b1c0_gen[22]),
                           .a23 (w_pr_pos_b1c0_gen[23]),
                           .a24 (w_pr_pos_b1c0_gen[24]),
                           .a25 (w_pr_pos_b1c0_gen[25]),
                           .a26 (w_pr_pos_b1c0_gen[26]),
                           .a27 (w_pr_pos_b1c0_gen[27]),
                           .a28 (w_pr_pos_b1c0_gen[28]),
                           .a29 (w_pr_pos_b1c0_gen[29]),
                           .a30 (w_pr_pos_b1c0_gen[30]),
                           .a31 (w_pr_pos_b1c0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_pos_b1c0));

//b1b0

generate
  for (i=0; i<32; i=i+1) begin : fetch_dec4
fetch_to_decode u_fetch_decode4 (.de_lower_16bytes  (        b1b0[((i*8)+31):i*8]), 
                                .w_pr_repne        (        w_pr_repne_b1b0_gen[i]),
                                .w_pr_cs_over      (      w_pr_cs_over_b1b0_gen[i]),
                                .w_pr_ss_over      (      w_pr_ss_over_b1b0_gen[i]),
                                .w_pr_ds_over      (      w_pr_ds_over_b1b0_gen[i]),
                                .w_pr_es_over      (      w_pr_es_over_b1b0_gen[i]),
                                .w_pr_fs_over      (      w_pr_fs_over_b1b0_gen[i]),
                                .w_pr_gs_over      (      w_pr_gs_over_b1b0_gen[i]),
                                .w_pr_size_over    (    w_pr_size_over_b1b0_gen[i]),
                                .w_pr_0f           (           w_pr_0f_b1b0_gen[i]),
                                .w_pr_pos          (          w_pr_pos_b1b0_gen[i]),
                                .w_mux_sel         (         w_mux_sel_b1b0_gen[i]));
  end
endgenerate

mux_nbit_32x1 #3 u_mux_sel4(.a0  (w_mux_sel_b1b0_gen[0 ]),  
                           .a1  (w_mux_sel_b1b0_gen[1 ]),
                           .a2  (w_mux_sel_b1b0_gen[2 ]),
                           .a3  (w_mux_sel_b1b0_gen[3 ]),
                           .a4  (w_mux_sel_b1b0_gen[4 ]),
                           .a5  (w_mux_sel_b1b0_gen[5 ]),
                           .a6  (w_mux_sel_b1b0_gen[6 ]),
                           .a7  (w_mux_sel_b1b0_gen[7 ]),
                           .a8  (w_mux_sel_b1b0_gen[8 ]),
                           .a9  (w_mux_sel_b1b0_gen[9 ]),
                           .a10 (w_mux_sel_b1b0_gen[10]),
                           .a11 (w_mux_sel_b1b0_gen[11]),
                           .a12 (w_mux_sel_b1b0_gen[12]),
                           .a13 (w_mux_sel_b1b0_gen[13]),
                           .a14 (w_mux_sel_b1b0_gen[14]),
                           .a15 (w_mux_sel_b1b0_gen[15]),
                           .a16 (w_mux_sel_b1b0_gen[16]),
                           .a17 (w_mux_sel_b1b0_gen[17]),
                           .a18 (w_mux_sel_b1b0_gen[18]),
                           .a19 (w_mux_sel_b1b0_gen[19]),
                           .a20 (w_mux_sel_b1b0_gen[20]),
                           .a21 (w_mux_sel_b1b0_gen[21]),
                           .a22 (w_mux_sel_b1b0_gen[22]),
                           .a23 (w_mux_sel_b1b0_gen[23]),
                           .a24 (w_mux_sel_b1b0_gen[24]),
                           .a25 (w_mux_sel_b1b0_gen[25]),
                           .a26 (w_mux_sel_b1b0_gen[26]),
                           .a27 (w_mux_sel_b1b0_gen[27]),
                           .a28 (w_mux_sel_b1b0_gen[28]),
                           .a29 (w_mux_sel_b1b0_gen[29]),
                           .a30 (w_mux_sel_b1b0_gen[30]),
                           .a31 (w_mux_sel_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_mux_sel_b1b0));


mux_nbit_32x1 #4 u_pr_repn4(.a0  (w_pr_repne_b1b0_gen[0 ]),  
                           .a1  (w_pr_repne_b1b0_gen[1 ]),
                           .a2  (w_pr_repne_b1b0_gen[2 ]),
                           .a3  (w_pr_repne_b1b0_gen[3 ]),
                           .a4  (w_pr_repne_b1b0_gen[4 ]),
                           .a5  (w_pr_repne_b1b0_gen[5 ]),
                           .a6  (w_pr_repne_b1b0_gen[6 ]),
                           .a7  (w_pr_repne_b1b0_gen[7 ]),
                           .a8  (w_pr_repne_b1b0_gen[8 ]),
                           .a9  (w_pr_repne_b1b0_gen[9 ]),
                           .a10 (w_pr_repne_b1b0_gen[10]),
                           .a11 (w_pr_repne_b1b0_gen[11]),
                           .a12 (w_pr_repne_b1b0_gen[12]),
                           .a13 (w_pr_repne_b1b0_gen[13]),
                           .a14 (w_pr_repne_b1b0_gen[14]),
                           .a15 (w_pr_repne_b1b0_gen[15]),
                           .a16 (w_pr_repne_b1b0_gen[16]),
                           .a17 (w_pr_repne_b1b0_gen[17]),
                           .a18 (w_pr_repne_b1b0_gen[18]),
                           .a19 (w_pr_repne_b1b0_gen[19]),
                           .a20 (w_pr_repne_b1b0_gen[20]),
                           .a21 (w_pr_repne_b1b0_gen[21]),
                           .a22 (w_pr_repne_b1b0_gen[22]),
                           .a23 (w_pr_repne_b1b0_gen[23]),
                           .a24 (w_pr_repne_b1b0_gen[24]),
                           .a25 (w_pr_repne_b1b0_gen[25]),
                           .a26 (w_pr_repne_b1b0_gen[26]),
                           .a27 (w_pr_repne_b1b0_gen[27]),
                           .a28 (w_pr_repne_b1b0_gen[28]),
                           .a29 (w_pr_repne_b1b0_gen[29]),
                           .a30 (w_pr_repne_b1b0_gen[30]),
                           .a31 (w_pr_repne_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_repne_b1b0));


mux_nbit_32x1 #4 u_pr_cs4  (.a0  (w_pr_cs_over_b1b0_gen[0 ]),  
                           .a1  (w_pr_cs_over_b1b0_gen[1 ]),
                           .a2  (w_pr_cs_over_b1b0_gen[2 ]),
                           .a3  (w_pr_cs_over_b1b0_gen[3 ]),
                           .a4  (w_pr_cs_over_b1b0_gen[4 ]),
                           .a5  (w_pr_cs_over_b1b0_gen[5 ]),
                           .a6  (w_pr_cs_over_b1b0_gen[6 ]),
                           .a7  (w_pr_cs_over_b1b0_gen[7 ]),
                           .a8  (w_pr_cs_over_b1b0_gen[8 ]),
                           .a9  (w_pr_cs_over_b1b0_gen[9 ]),
                           .a10 (w_pr_cs_over_b1b0_gen[10]),
                           .a11 (w_pr_cs_over_b1b0_gen[11]),
                           .a12 (w_pr_cs_over_b1b0_gen[12]),
                           .a13 (w_pr_cs_over_b1b0_gen[13]),
                           .a14 (w_pr_cs_over_b1b0_gen[14]),
                           .a15 (w_pr_cs_over_b1b0_gen[15]),
                           .a16 (w_pr_cs_over_b1b0_gen[16]),
                           .a17 (w_pr_cs_over_b1b0_gen[17]),
                           .a18 (w_pr_cs_over_b1b0_gen[18]),
                           .a19 (w_pr_cs_over_b1b0_gen[19]),
                           .a20 (w_pr_cs_over_b1b0_gen[20]),
                           .a21 (w_pr_cs_over_b1b0_gen[21]),
                           .a22 (w_pr_cs_over_b1b0_gen[22]),
                           .a23 (w_pr_cs_over_b1b0_gen[23]),
                           .a24 (w_pr_cs_over_b1b0_gen[24]),
                           .a25 (w_pr_cs_over_b1b0_gen[25]),
                           .a26 (w_pr_cs_over_b1b0_gen[26]),
                           .a27 (w_pr_cs_over_b1b0_gen[27]),
                           .a28 (w_pr_cs_over_b1b0_gen[28]),
                           .a29 (w_pr_cs_over_b1b0_gen[29]),
                           .a30 (w_pr_cs_over_b1b0_gen[30]),
                           .a31 (w_pr_cs_over_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_cs_over_b1b0));

mux_nbit_32x1 #4 u_pr_ss4  (.a0  (w_pr_ss_over_b1b0_gen[0 ]),  
                           .a1  (w_pr_ss_over_b1b0_gen[1 ]),
                           .a2  (w_pr_ss_over_b1b0_gen[2 ]),
                           .a3  (w_pr_ss_over_b1b0_gen[3 ]),
                           .a4  (w_pr_ss_over_b1b0_gen[4 ]),
                           .a5  (w_pr_ss_over_b1b0_gen[5 ]),
                           .a6  (w_pr_ss_over_b1b0_gen[6 ]),
                           .a7  (w_pr_ss_over_b1b0_gen[7 ]),
                           .a8  (w_pr_ss_over_b1b0_gen[8 ]),
                           .a9  (w_pr_ss_over_b1b0_gen[9 ]),
                           .a10 (w_pr_ss_over_b1b0_gen[10]),
                           .a11 (w_pr_ss_over_b1b0_gen[11]),
                           .a12 (w_pr_ss_over_b1b0_gen[12]),
                           .a13 (w_pr_ss_over_b1b0_gen[13]),
                           .a14 (w_pr_ss_over_b1b0_gen[14]),
                           .a15 (w_pr_ss_over_b1b0_gen[15]),
                           .a16 (w_pr_ss_over_b1b0_gen[16]),
                           .a17 (w_pr_ss_over_b1b0_gen[17]),
                           .a18 (w_pr_ss_over_b1b0_gen[18]),
                           .a19 (w_pr_ss_over_b1b0_gen[19]),
                           .a20 (w_pr_ss_over_b1b0_gen[20]),
                           .a21 (w_pr_ss_over_b1b0_gen[21]),
                           .a22 (w_pr_ss_over_b1b0_gen[22]),
                           .a23 (w_pr_ss_over_b1b0_gen[23]),
                           .a24 (w_pr_ss_over_b1b0_gen[24]),
                           .a25 (w_pr_ss_over_b1b0_gen[25]),
                           .a26 (w_pr_ss_over_b1b0_gen[26]),
                           .a27 (w_pr_ss_over_b1b0_gen[27]),
                           .a28 (w_pr_ss_over_b1b0_gen[28]),
                           .a29 (w_pr_ss_over_b1b0_gen[29]),
                           .a30 (w_pr_ss_over_b1b0_gen[30]),
                           .a31 (w_pr_ss_over_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ss_over_b1b0));

mux_nbit_32x1 #4 u_pr_ds4  (.a0  (w_pr_ds_over_b1b0_gen[0 ]),  
                           .a1  (w_pr_ds_over_b1b0_gen[1 ]),
                           .a2  (w_pr_ds_over_b1b0_gen[2 ]),
                           .a3  (w_pr_ds_over_b1b0_gen[3 ]),
                           .a4  (w_pr_ds_over_b1b0_gen[4 ]),
                           .a5  (w_pr_ds_over_b1b0_gen[5 ]),
                           .a6  (w_pr_ds_over_b1b0_gen[6 ]),
                           .a7  (w_pr_ds_over_b1b0_gen[7 ]),
                           .a8  (w_pr_ds_over_b1b0_gen[8 ]),
                           .a9  (w_pr_ds_over_b1b0_gen[9 ]),
                           .a10 (w_pr_ds_over_b1b0_gen[10]),
                           .a11 (w_pr_ds_over_b1b0_gen[11]),
                           .a12 (w_pr_ds_over_b1b0_gen[12]),
                           .a13 (w_pr_ds_over_b1b0_gen[13]),
                           .a14 (w_pr_ds_over_b1b0_gen[14]),
                           .a15 (w_pr_ds_over_b1b0_gen[15]),
                           .a16 (w_pr_ds_over_b1b0_gen[16]),
                           .a17 (w_pr_ds_over_b1b0_gen[17]),
                           .a18 (w_pr_ds_over_b1b0_gen[18]),
                           .a19 (w_pr_ds_over_b1b0_gen[19]),
                           .a20 (w_pr_ds_over_b1b0_gen[20]),
                           .a21 (w_pr_ds_over_b1b0_gen[21]),
                           .a22 (w_pr_ds_over_b1b0_gen[22]),
                           .a23 (w_pr_ds_over_b1b0_gen[23]),
                           .a24 (w_pr_ds_over_b1b0_gen[24]),
                           .a25 (w_pr_ds_over_b1b0_gen[25]),
                           .a26 (w_pr_ds_over_b1b0_gen[26]),
                           .a27 (w_pr_ds_over_b1b0_gen[27]),
                           .a28 (w_pr_ds_over_b1b0_gen[28]),
                           .a29 (w_pr_ds_over_b1b0_gen[29]),
                           .a30 (w_pr_ds_over_b1b0_gen[30]),
                           .a31 (w_pr_ds_over_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_ds_over_b1b0));

mux_nbit_32x1 #4 u_pr_es4  (.a0  (w_pr_es_over_b1b0_gen[0 ]),  
                           .a1  (w_pr_es_over_b1b0_gen[1 ]),
                           .a2  (w_pr_es_over_b1b0_gen[2 ]),
                           .a3  (w_pr_es_over_b1b0_gen[3 ]),
                           .a4  (w_pr_es_over_b1b0_gen[4 ]),
                           .a5  (w_pr_es_over_b1b0_gen[5 ]),
                           .a6  (w_pr_es_over_b1b0_gen[6 ]),
                           .a7  (w_pr_es_over_b1b0_gen[7 ]),
                           .a8  (w_pr_es_over_b1b0_gen[8 ]),
                           .a9  (w_pr_es_over_b1b0_gen[9 ]),
                           .a10 (w_pr_es_over_b1b0_gen[10]),
                           .a11 (w_pr_es_over_b1b0_gen[11]),
                           .a12 (w_pr_es_over_b1b0_gen[12]),
                           .a13 (w_pr_es_over_b1b0_gen[13]),
                           .a14 (w_pr_es_over_b1b0_gen[14]),
                           .a15 (w_pr_es_over_b1b0_gen[15]),
                           .a16 (w_pr_es_over_b1b0_gen[16]),
                           .a17 (w_pr_es_over_b1b0_gen[17]),
                           .a18 (w_pr_es_over_b1b0_gen[18]),
                           .a19 (w_pr_es_over_b1b0_gen[19]),
                           .a20 (w_pr_es_over_b1b0_gen[20]),
                           .a21 (w_pr_es_over_b1b0_gen[21]),
                           .a22 (w_pr_es_over_b1b0_gen[22]),
                           .a23 (w_pr_es_over_b1b0_gen[23]),
                           .a24 (w_pr_es_over_b1b0_gen[24]),
                           .a25 (w_pr_es_over_b1b0_gen[25]),
                           .a26 (w_pr_es_over_b1b0_gen[26]),
                           .a27 (w_pr_es_over_b1b0_gen[27]),
                           .a28 (w_pr_es_over_b1b0_gen[28]),
                           .a29 (w_pr_es_over_b1b0_gen[29]),
                           .a30 (w_pr_es_over_b1b0_gen[30]),
                           .a31 (w_pr_es_over_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_es_over_b1b0));

mux_nbit_32x1 #4 u_pr_fs4  (.a0  (w_pr_fs_over_b1b0_gen[0 ]),  
                           .a1  (w_pr_fs_over_b1b0_gen[1 ]),
                           .a2  (w_pr_fs_over_b1b0_gen[2 ]),
                           .a3  (w_pr_fs_over_b1b0_gen[3 ]),
                           .a4  (w_pr_fs_over_b1b0_gen[4 ]),
                           .a5  (w_pr_fs_over_b1b0_gen[5 ]),
                           .a6  (w_pr_fs_over_b1b0_gen[6 ]),
                           .a7  (w_pr_fs_over_b1b0_gen[7 ]),
                           .a8  (w_pr_fs_over_b1b0_gen[8 ]),
                           .a9  (w_pr_fs_over_b1b0_gen[9 ]),
                           .a10 (w_pr_fs_over_b1b0_gen[10]),
                           .a11 (w_pr_fs_over_b1b0_gen[11]),
                           .a12 (w_pr_fs_over_b1b0_gen[12]),
                           .a13 (w_pr_fs_over_b1b0_gen[13]),
                           .a14 (w_pr_fs_over_b1b0_gen[14]),
                           .a15 (w_pr_fs_over_b1b0_gen[15]),
                           .a16 (w_pr_fs_over_b1b0_gen[16]),
                           .a17 (w_pr_fs_over_b1b0_gen[17]),
                           .a18 (w_pr_fs_over_b1b0_gen[18]),
                           .a19 (w_pr_fs_over_b1b0_gen[19]),
                           .a20 (w_pr_fs_over_b1b0_gen[20]),
                           .a21 (w_pr_fs_over_b1b0_gen[21]),
                           .a22 (w_pr_fs_over_b1b0_gen[22]),
                           .a23 (w_pr_fs_over_b1b0_gen[23]),
                           .a24 (w_pr_fs_over_b1b0_gen[24]),
                           .a25 (w_pr_fs_over_b1b0_gen[25]),
                           .a26 (w_pr_fs_over_b1b0_gen[26]),
                           .a27 (w_pr_fs_over_b1b0_gen[27]),
                           .a28 (w_pr_fs_over_b1b0_gen[28]),
                           .a29 (w_pr_fs_over_b1b0_gen[29]),
                           .a30 (w_pr_fs_over_b1b0_gen[30]),
                           .a31 (w_pr_fs_over_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_fs_over_b1b0));

mux_nbit_32x1 #4 u_pr_gs4  (.a0  (w_pr_gs_over_b1b0_gen[0 ]),  
                           .a1  (w_pr_gs_over_b1b0_gen[1 ]),
                           .a2  (w_pr_gs_over_b1b0_gen[2 ]),
                           .a3  (w_pr_gs_over_b1b0_gen[3 ]),
                           .a4  (w_pr_gs_over_b1b0_gen[4 ]),
                           .a5  (w_pr_gs_over_b1b0_gen[5 ]),
                           .a6  (w_pr_gs_over_b1b0_gen[6 ]),
                           .a7  (w_pr_gs_over_b1b0_gen[7 ]),
                           .a8  (w_pr_gs_over_b1b0_gen[8 ]),
                           .a9  (w_pr_gs_over_b1b0_gen[9 ]),
                           .a10 (w_pr_gs_over_b1b0_gen[10]),
                           .a11 (w_pr_gs_over_b1b0_gen[11]),
                           .a12 (w_pr_gs_over_b1b0_gen[12]),
                           .a13 (w_pr_gs_over_b1b0_gen[13]),
                           .a14 (w_pr_gs_over_b1b0_gen[14]),
                           .a15 (w_pr_gs_over_b1b0_gen[15]),
                           .a16 (w_pr_gs_over_b1b0_gen[16]),
                           .a17 (w_pr_gs_over_b1b0_gen[17]),
                           .a18 (w_pr_gs_over_b1b0_gen[18]),
                           .a19 (w_pr_gs_over_b1b0_gen[19]),
                           .a20 (w_pr_gs_over_b1b0_gen[20]),
                           .a21 (w_pr_gs_over_b1b0_gen[21]),
                           .a22 (w_pr_gs_over_b1b0_gen[22]),
                           .a23 (w_pr_gs_over_b1b0_gen[23]),
                           .a24 (w_pr_gs_over_b1b0_gen[24]),
                           .a25 (w_pr_gs_over_b1b0_gen[25]),
                           .a26 (w_pr_gs_over_b1b0_gen[26]),
                           .a27 (w_pr_gs_over_b1b0_gen[27]),
                           .a28 (w_pr_gs_over_b1b0_gen[28]),
                           .a29 (w_pr_gs_over_b1b0_gen[29]),
                           .a30 (w_pr_gs_over_b1b0_gen[30]),
                           .a31 (w_pr_gs_over_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_gs_over_b1b0));

mux_nbit_32x1 #4 u_pr_size4(.a0  (w_pr_size_over_b1b0_gen[0 ]),  
                           .a1  (w_pr_size_over_b1b0_gen[1 ]),
                           .a2  (w_pr_size_over_b1b0_gen[2 ]),
                           .a3  (w_pr_size_over_b1b0_gen[3 ]),
                           .a4  (w_pr_size_over_b1b0_gen[4 ]),
                           .a5  (w_pr_size_over_b1b0_gen[5 ]),
                           .a6  (w_pr_size_over_b1b0_gen[6 ]),
                           .a7  (w_pr_size_over_b1b0_gen[7 ]),
                           .a8  (w_pr_size_over_b1b0_gen[8 ]),
                           .a9  (w_pr_size_over_b1b0_gen[9 ]),
                           .a10 (w_pr_size_over_b1b0_gen[10]),
                           .a11 (w_pr_size_over_b1b0_gen[11]),
                           .a12 (w_pr_size_over_b1b0_gen[12]),
                           .a13 (w_pr_size_over_b1b0_gen[13]),
                           .a14 (w_pr_size_over_b1b0_gen[14]),
                           .a15 (w_pr_size_over_b1b0_gen[15]),
                           .a16 (w_pr_size_over_b1b0_gen[16]),
                           .a17 (w_pr_size_over_b1b0_gen[17]),
                           .a18 (w_pr_size_over_b1b0_gen[18]),
                           .a19 (w_pr_size_over_b1b0_gen[19]),
                           .a20 (w_pr_size_over_b1b0_gen[20]),
                           .a21 (w_pr_size_over_b1b0_gen[21]),
                           .a22 (w_pr_size_over_b1b0_gen[22]),
                           .a23 (w_pr_size_over_b1b0_gen[23]),
                           .a24 (w_pr_size_over_b1b0_gen[24]),
                           .a25 (w_pr_size_over_b1b0_gen[25]),
                           .a26 (w_pr_size_over_b1b0_gen[26]),
                           .a27 (w_pr_size_over_b1b0_gen[27]),
                           .a28 (w_pr_size_over_b1b0_gen[28]),
                           .a29 (w_pr_size_over_b1b0_gen[29]),
                           .a30 (w_pr_size_over_b1b0_gen[30]),
                           .a31 (w_pr_size_over_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_size_over_b1b0));

mux_nbit_32x1 #4 u_pr_0f4  (.a0  (w_pr_0f_b1b0_gen[0 ]),  
                           .a1  (w_pr_0f_b1b0_gen[1 ]),
                           .a2  (w_pr_0f_b1b0_gen[2 ]),
                           .a3  (w_pr_0f_b1b0_gen[3 ]),
                           .a4  (w_pr_0f_b1b0_gen[4 ]),
                           .a5  (w_pr_0f_b1b0_gen[5 ]),
                           .a6  (w_pr_0f_b1b0_gen[6 ]),
                           .a7  (w_pr_0f_b1b0_gen[7 ]),
                           .a8  (w_pr_0f_b1b0_gen[8 ]),
                           .a9  (w_pr_0f_b1b0_gen[9 ]),
                           .a10 (w_pr_0f_b1b0_gen[10]),
                           .a11 (w_pr_0f_b1b0_gen[11]),
                           .a12 (w_pr_0f_b1b0_gen[12]),
                           .a13 (w_pr_0f_b1b0_gen[13]),
                           .a14 (w_pr_0f_b1b0_gen[14]),
                           .a15 (w_pr_0f_b1b0_gen[15]),
                           .a16 (w_pr_0f_b1b0_gen[16]),
                           .a17 (w_pr_0f_b1b0_gen[17]),
                           .a18 (w_pr_0f_b1b0_gen[18]),
                           .a19 (w_pr_0f_b1b0_gen[19]),
                           .a20 (w_pr_0f_b1b0_gen[20]),
                           .a21 (w_pr_0f_b1b0_gen[21]),
                           .a22 (w_pr_0f_b1b0_gen[22]),
                           .a23 (w_pr_0f_b1b0_gen[23]),
                           .a24 (w_pr_0f_b1b0_gen[24]),
                           .a25 (w_pr_0f_b1b0_gen[25]),
                           .a26 (w_pr_0f_b1b0_gen[26]),
                           .a27 (w_pr_0f_b1b0_gen[27]),
                           .a28 (w_pr_0f_b1b0_gen[28]),
                           .a29 (w_pr_0f_b1b0_gen[29]),
                           .a30 (w_pr_0f_b1b0_gen[30]),
                           .a31 (w_pr_0f_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_0f_b1b0));

mux_nbit_32x1 #4 u_pr_pos4 (.a0  (w_pr_pos_b1b0_gen[0 ]),  
                           .a1  (w_pr_pos_b1b0_gen[1 ]),
                           .a2  (w_pr_pos_b1b0_gen[2 ]),
                           .a3  (w_pr_pos_b1b0_gen[3 ]),
                           .a4  (w_pr_pos_b1b0_gen[4 ]),
                           .a5  (w_pr_pos_b1b0_gen[5 ]),
                           .a6  (w_pr_pos_b1b0_gen[6 ]),
                           .a7  (w_pr_pos_b1b0_gen[7 ]),
                           .a8  (w_pr_pos_b1b0_gen[8 ]),
                           .a9  (w_pr_pos_b1b0_gen[9 ]),
                           .a10 (w_pr_pos_b1b0_gen[10]),
                           .a11 (w_pr_pos_b1b0_gen[11]),
                           .a12 (w_pr_pos_b1b0_gen[12]),
                           .a13 (w_pr_pos_b1b0_gen[13]),
                           .a14 (w_pr_pos_b1b0_gen[14]),
                           .a15 (w_pr_pos_b1b0_gen[15]),
                           .a16 (w_pr_pos_b1b0_gen[16]),
                           .a17 (w_pr_pos_b1b0_gen[17]),
                           .a18 (w_pr_pos_b1b0_gen[18]),
                           .a19 (w_pr_pos_b1b0_gen[19]),
                           .a20 (w_pr_pos_b1b0_gen[20]),
                           .a21 (w_pr_pos_b1b0_gen[21]),
                           .a22 (w_pr_pos_b1b0_gen[22]),
                           .a23 (w_pr_pos_b1b0_gen[23]),
                           .a24 (w_pr_pos_b1b0_gen[24]),
                           .a25 (w_pr_pos_b1b0_gen[25]),
                           .a26 (w_pr_pos_b1b0_gen[26]),
                           .a27 (w_pr_pos_b1b0_gen[27]),
                           .a28 (w_pr_pos_b1b0_gen[28]),
                           .a29 (w_pr_pos_b1b0_gen[29]),
                           .a30 (w_pr_pos_b1b0_gen[30]),
                           .a31 (w_pr_pos_b1b0_gen[31]),
                           .sel (w_EIP_to_use[4:0]),
                           .out (w_pr_pos_b1b0));


mux_nbit_4x1 #3 u_1(.a0(w_mux_sel_b1b0), .a1(w_mux_sel_b1c0), .a2(w_mux_sel_c1b0), .a3(w_mux_sel_c1c0), .sel(w_fe_ld_buf), .out(w_mux_sel));

mux_nbit_4x1 #4 u_2(.a0(w_pr_repne_b1b0), .a1(w_pr_repne_b1c0), .a2(w_pr_repne_c1b0), .a3(w_pr_repne_c1c0), .sel(w_fe_ld_buf), .out(w_pr_repne));

mux_nbit_4x1 #4 u_3(.a0(w_pr_cs_over_b1b0), .a1(w_pr_cs_over_b1c0), .a2(w_pr_cs_over_c1b0), .a3(w_pr_cs_over_c1c0), .sel(w_fe_ld_buf), .out(w_pr_cs_over));

mux_nbit_4x1 #4 u_4(.a0(w_pr_ss_over_b1b0), .a1(w_pr_ss_over_b1c0), .a2(w_pr_ss_over_c1b0), .a3(w_pr_ss_over_c1c0), .sel(w_fe_ld_buf), .out(w_pr_ss_over));

mux_nbit_4x1 #4 u_5(.a0(w_pr_ds_over_b1b0), .a1(w_pr_ds_over_b1c0), .a2(w_pr_ds_over_c1b0), .a3(w_pr_ds_over_c1c0), .sel(w_fe_ld_buf), .out(w_pr_ds_over));

mux_nbit_4x1 #4 u_6(.a0(w_pr_es_over_b1b0), .a1(w_pr_es_over_b1c0), .a2(w_pr_es_over_c1b0), .a3(w_pr_es_over_c1c0), .sel(w_fe_ld_buf), .out(w_pr_es_over));

mux_nbit_4x1 #4 u_7(.a0(w_pr_fs_over_b1b0), .a1(w_pr_fs_over_b1c0), .a2(w_pr_fs_over_c1b0), .a3(w_pr_fs_over_c1c0), .sel(w_fe_ld_buf), .out(w_pr_fs_over));

mux_nbit_4x1 #4 u_8(.a0(w_pr_gs_over_b1b0), .a1(w_pr_gs_over_b1c0), .a2(w_pr_gs_over_c1b0), .a3(w_pr_gs_over_c1c0), .sel(w_fe_ld_buf), .out(w_pr_gs_over));

mux_nbit_4x1 #4 u_9(.a0(w_pr_size_over_b1b0), .a1(w_pr_size_over_b1c0), .a2(w_pr_size_over_c1b0), .a3(w_pr_size_over_c1c0), .sel(w_fe_ld_buf), .out(w_pr_size_over));

mux_nbit_4x1 #4 u_10(.a0(w_pr_0f_b1b0), .a1(w_pr_0f_b1c0), .a2(w_pr_0f_c1b0), .a3(w_pr_0f_c1c0), .sel(w_fe_ld_buf), .out(w_pr_0f));

mux_nbit_4x1 #4 u_11(.a0(w_pr_pos_b1b0), .a1(w_pr_pos_b1c0), .a2(w_pr_pos_c1b0), .a3(w_pr_pos_c1c0), .sel(w_fe_ld_buf), .out(w_pr_pos));

endmodule
