module cpu_top
(
  input clk,
  input rst_n
);

// ********** Hardcoded entries ***********
//TLB entries
reg [7:0] TLB[31:0]; //actually 30 bit entries

//Segment_limit_Regs
reg [31:0] CS_limit;

initial begin
  TLB[0] = 32'h0000;
  TLB[1] = 32'h0000;
  TLB[2] = 32'h0000;
  TLB[3] = 32'h0000;
  TLB[4] = 32'h0000;
  TLB[5] = 32'h0000;
  TLB[6] = 32'h0000;
  TLB[7] = 32'h0000;
  
  CS_limit = 32'h3ff;
end


//Signals between fetch and decode
//Output of fetch
wire [127:0] de_lower_data;
wire [127:0] de_upper_data;

//Input to fetch
wire de_p;

wire [31:0] wb_data1;

// ***************** FETCH STAGE ******************

wire EIP_1, not_EIP_1;
wire [1:0] f_state;
wire [31:0] f_address;
wire [2:0] f_PFN;
wire [1:0] f_ld_buf;
wire [127:0] icache_lower_data;
wire [127:0] icache_upper_data;
wire [127:0] icache_lower_data_reg;
wire [127:0] icache_upper_data_reg;
wire [127:0] icache_shifted_lower_data;
wire [127:0] icache_shifted_upper_data;

// EIP register
wire ld_EIP;
wire [31:0] EIP_reg;
wire [31:0] EIP_updated;
wire [31:0] next_EIP;
wire EIP_mux;
register u_EIP(clk, rst_n, 1'b1, EIP_updated, EIP_reg, ld_EIP);
mux_nbit_2x1 #32 u_EIP_updated (next_EIP, wb_data1, EIP_mux, EIP_updated);

wire [31:0] EIP_plus_32;
kogge_stone #32 u_EIP_reg (EIP_reg, 32'h10, 1'b0, EIP_plus_32, , ); 

// 2nd register
wire f_second_updated;
wire f_second_reg;
wire f_second_int; //Generated by fetch fsm
NOT u_not_f_second_reg (f_second_reg, not_f_second_reg);
nor2$ u_state_is_00 (state_is_00, f_state[0], f_state[1]);
and2$ u_f_second_int (f_second_int, state_is_00, EIP_1);

and2$ u_f_second_updated (f_second_updated, not_f_second_reg, f_second_int);
register #1 u_f_second_reg (clk, rst_n, 1'b1, f_second_updated, f_second_reg, 1'b1);

//EIP_1
assign EIP_1 = EIP_reg[4];

// fetch_address
wire f_address_sel; // (state==00 && (!eip_1 || f_second_updated))
wire w_eip0_or_second;
or2$ u_w_eip0_or_second (w_eip0_or_second, not_EIP_1, f_second_updated);
and2$ u_f_address_sel (f_address_sel, w_eip0_or_second, state_is_00);
mux_nbit_2x1 #32 u_f_address( EIP_plus_32, EIP_reg, f_address_sel, f_address);

//ren //FIXME: not of all future stalls and not int_trig
assign f_ren = 1'b1; 

// Fetch FSM
fetch_fsm u_fetch_fsm (
  .clk      (clk),
  .rst_n    (rst_n),
  .second   (f_second_updated),
  .de_p     (de_p),
  .eip_4    (EIP_reg[4]),
  .ld_buf   (f_ld_buf),
  .curr_st  (f_state)
  );

//Instruction cache
i_cache u_i_cache (
  .clk          (clk),
  .ren          (f_ren),
  .index        (f_address[8:5]),
  .tag_14_12    (f_PFN),
  .tag_11_9     (f_address[11:9]),
  .ic_fill_data (),
  .ic_miss_ack  (),
  .v_init       (),
  .r_data       (),
  .r_ready      (),
  .ic_miss      (),
  .ic_addr      ()
);              

//Logic that checks TLB entries and gives the PFN, exceptions
wire [7:0] f_TLB_hits;
wire f_TLB_hit;
genvar i;
generate begin : loop
for (i=0; i<8; i=i+1) begin
  eq_checker #25 ({TLB[i][29:7], TLB[i][4], TLB[i][3]}, {f_address[31:9],1'b1,1'b1}, f_TLB_hits[i]);
end
end
endgenerate

wire in_CS_limit;
//FIXME : need to write <, > submodules
assign in_CS_limit = (f_address < CS_limit);
wire in_CS_limit_and_ren;
and2$ u_in_CS_limit_and_ren( in_CS_limit_and_ren, in_CS_limit, f_ren);

wire [1:0] w_f_tlbhit;
and4$ u_w_tlbhit0 (w_f_tlbhit[0], f_TLB_hits[0], f_TLB_hits[1], f_TLB_hits[2], f_TLB_hits[3]);
and4$ u_w_tlbhit1 (w_f_tlbhit[1], f_TLB_hits[4], f_TLB_hits[5], f_TLB_hits[6], f_TLB_hits[7]);
and2$ u_f_TLB_hit (f_TLB_hit, w_f_tlbhit[0], w_f_tlbhit[1]);

wire f_pg_fault;
and2$ u_f_pg_fault (f_pg_fault, in_CS_limit_and_ren, f_TLB_hit);

mux_nbit_8x1_mulsel #3 u_f_pfn (TLB[0][6:4], TLB[1][6:4], TLB[2][6:4], TLB[3][6:4], 
                        TLB[4][6:4], TLB[5][6:4], TLB[6][6:4], TLB[7][6:4], 
                        f_TLB_hits[0], f_TLB_hits[1], f_TLB_hits[2], f_TLB_hits[3], 
                        f_TLB_hits[4], f_TLB_hits[5], f_TLB_hits[6], f_TLB_hits[7], f_PFN);


//Latching icache data
register #128 u_i_lower_data_reg (clk, rst_n, 1'b1, icache_lower_data, icache_lower_data_reg, f_ld_buf[0]);
register #128 u_i_upper_data_reg (clk, rst_n, 1'b1, icache_upper_data, icache_upper_data_reg, f_ld_buf[1]);

//shifted icache data
//FIXME : need to multiply EIP with 8, and need shift right rotate
shift_right #256 u_i_shifter_ldata (
  .amt(EIP_reg[4:0]),
  .sin(1'b0),
  .in({icache_upper_data, icache_lower_data}),
  .out({icache_shifted_upper_data, icache_shifted_lower_data}),
  .sout()
  );


// ***************** WRITEBACK STAGE ******************


endmodule


